* File: ROM_MACRO.pex.spi
* Created: Mon Jan 17 05:42:50 2022
* Program "Calibre xRC"
* Version "v2021.1_33.19"
* 
.include "ROM_MACRO.pex.spi.pex"
.subckt ROM_MACRO  VSS CLK VDD VREF A<7> A<6> A<2> A<1> A<0> DOUT<1> A<8> A<5>
+ A<4> A<3> DOUT<0>
* 
* DOUT<0>	DOUT<0>
* A<3>	A<3>
* A<4>	A<4>
* A<5>	A<5>
* A<8>	A<8>
* DOUT<1>	DOUT<1>
* A<0>	A<0>
* A<1>	A<1>
* A<2>	A<2>
* A<6>	A<6>
* A<7>	A<7>
* VREF	VREF
* VDD	VDD
* CLK	CLK
* VSS	VSS
mXI45/XI0/XI8/MM0 N_XI45/XI0/NET96_XI45/XI0/XI8/MM0_d
+ N_NET100_XI45/XI0/XI8/MM0_g N_VSS_XI45/XI0/XI8/MM0_s N_VSS_XI45/XI0/XI8/MM0_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI45/XI1/XI8/MM0 N_XI45/XI1/NET96_XI45/XI1/XI8/MM0_d
+ N_NET110_XI45/XI1/XI8/MM0_g N_VSS_XI45/XI1/XI8/MM0_s N_VSS_XI45/XI0/XI8/MM0_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI46/MM3 N_NET0208_XI46/MM3_d N_NET0265_XI46/MM3_g N_DOUT<1>_XI46/MM3_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=7.5e-07 AD=3.675e-13 AS=1.92e-13
+ PD=1.73e-06 PS=8.58e-07
mXI46/MM1 N_DOUT<1>_XI46/MM1_d N_NET0176_XI46/MM1_g N_VSS_XI46/MM1_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.28e-13 AS=1.8e-13
+ PD=5.72e-07 PS=7.2e-07
mXI46/MM2 N_NET0176_XI46/MM2_d N_DOUT<1>_XI46/MM2_g N_VSS_XI46/MM2_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.28e-13 AS=1.8e-13
+ PD=5.72e-07 PS=7.2e-07
mXI46/MM0 N_NET0207_XI46/MM0_d N_NET0265_XI46/MM0_g N_NET0176_XI46/MM0_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=7.5e-07 AD=3.675e-13 AS=1.92e-13
+ PD=1.73e-06 PS=8.58e-07
mXI10/MM7 N_XI10/NET13_XI10/MM7_d N_A<7>_XI10/MM7_g N_VSS_XI10/MM7_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI10/MM8 N_XI10/NET9_XI10/MM8_d N_CLK_XI10/MM8_g N_VSS_XI10/MM8_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI10/MM5 N_XI10/NET21_XI10/MM5_d N_XI10/NET13_XI10/MM5_g N_XI10/NET9_XI10/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI10/MM9 N_XI10/NET5_XI10/MM9_d N_XI10/NET21_XI10/MM9_g N_VSS_XI10/MM9_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI10/MM6 N_XI10/NET15_XI10/MM6_d N_CLK_XI10/MM6_g N_XI10/NET5_XI10/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI10/MM10 N_NET125_XI10/MM10_d N_XI10/NET15_XI10/MM10_g N_VSS_XI10/MM10_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI18/MM7 N_XI18/NET13_XI18/MM7_d N_A<6>_XI18/MM7_g N_VSS_XI18/MM7_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI18/MM8 N_XI18/NET9_XI18/MM8_d N_CLK_XI18/MM8_g N_VSS_XI18/MM8_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI18/MM5 N_XI18/NET21_XI18/MM5_d N_XI18/NET13_XI18/MM5_g N_XI18/NET9_XI18/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI18/MM9 N_XI18/NET5_XI18/MM9_d N_XI18/NET21_XI18/MM9_g N_VSS_XI18/MM9_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI18/MM6 N_XI18/NET15_XI18/MM6_d N_CLK_XI18/MM6_g N_XI18/NET5_XI18/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI18/MM10 N_NET85_XI18/MM10_d N_XI18/NET15_XI18/MM10_g N_VSS_XI18/MM10_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI16/MM7 N_XI16/NET13_XI16/MM7_d N_A<2>_XI16/MM7_g N_VSS_XI16/MM7_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI16/MM8 N_XI16/NET9_XI16/MM8_d N_CLK_XI16/MM8_g N_VSS_XI16/MM8_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI16/MM5 N_XI16/NET21_XI16/MM5_d N_XI16/NET13_XI16/MM5_g N_XI16/NET9_XI16/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI16/MM9 N_XI16/NET5_XI16/MM9_d N_XI16/NET21_XI16/MM9_g N_VSS_XI16/MM9_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI16/MM6 N_XI16/NET15_XI16/MM6_d N_CLK_XI16/MM6_g N_XI16/NET5_XI16/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI16/MM10 N_NET95_XI16/MM10_d N_XI16/NET15_XI16/MM10_g N_VSS_XI16/MM10_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI14/MM7 N_XI14/NET13_XI14/MM7_d N_A<1>_XI14/MM7_g N_VSS_XI14/MM7_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI14/MM8 N_XI14/NET9_XI14/MM8_d N_CLK_XI14/MM8_g N_VSS_XI14/MM8_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI14/MM5 N_XI14/NET21_XI14/MM5_d N_XI14/NET13_XI14/MM5_g N_XI14/NET9_XI14/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI14/MM9 N_XI14/NET5_XI14/MM9_d N_XI14/NET21_XI14/MM9_g N_VSS_XI14/MM9_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI14/MM6 N_XI14/NET15_XI14/MM6_d N_CLK_XI14/MM6_g N_XI14/NET5_XI14/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI14/MM10 N_NET105_XI14/MM10_d N_XI14/NET15_XI14/MM10_g N_VSS_XI14/MM10_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI15/MM7 N_XI15/NET13_XI15/MM7_d N_A<0>_XI15/MM7_g N_VSS_XI15/MM7_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI15/MM8 N_XI15/NET9_XI15/MM8_d N_CLK_XI15/MM8_g N_VSS_XI15/MM8_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI15/MM5 N_XI15/NET21_XI15/MM5_d N_XI15/NET13_XI15/MM5_g N_XI15/NET9_XI15/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI15/MM9 N_XI15/NET5_XI15/MM9_d N_XI15/NET21_XI15/MM9_g N_VSS_XI15/MM9_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI15/MM6 N_XI15/NET15_XI15/MM6_d N_CLK_XI15/MM6_g N_XI15/NET5_XI15/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI15/MM10 N_NET100_XI15/MM10_d N_XI15/NET15_XI15/MM10_g N_VSS_XI15/MM10_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI45/XI0/XI9/MM0 N_XI45/XI0/NET92_XI45/XI0/XI9/MM0_d
+ N_NET105_XI45/XI0/XI9/MM0_g N_VSS_XI45/XI0/XI9/MM0_s N_VSS_XI45/XI0/XI8/MM0_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI45/XI1/XI9/MM0 N_XI45/XI1/NET92_XI45/XI1/XI9/MM0_d N_NET90_XI45/XI1/XI9/MM0_g
+ N_VSS_XI45/XI1/XI9/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI45/XI0/XI10/MM0 N_XI45/XI0/NET081_XI45/XI0/XI10/MM0_d
+ N_NET95_XI45/XI0/XI10/MM0_g N_VSS_XI45/XI0/XI10/MM0_s N_VSS_XI45/XI0/XI8/MM0_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI45/XI1/XI10/MM0 N_XI45/XI1/NET081_XI45/XI1/XI10/MM0_d
+ N_NET115_XI45/XI1/XI10/MM0_g N_VSS_XI45/XI1/XI10/MM0_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI45/XI0/XI18/MM7 N_XI45/NET272_XI45/XI0/XI18/MM7_d N_NET79_XI45/XI0/XI18/MM7_g
+ N_XI45/XI0/XI18/NET16_XI45/XI0/XI18/MM7_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI18/MM6 N_XI45/XI0/XI18/NET16_XI45/XI0/XI18/MM6_d
+ N_XI45/XI0/NET081_XI45/XI0/XI18/MM6_g
+ N_XI45/XI0/XI18/NET12_XI45/XI0/XI18/MM6_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI18/MM5 N_XI45/XI0/XI18/NET12_XI45/XI0/XI18/MM5_d
+ N_XI45/XI0/NET92_XI45/XI0/XI18/MM5_g N_XI45/XI0/XI18/NET8_XI45/XI0/XI18/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI18/MM4 N_XI45/XI0/XI18/NET8_XI45/XI0/XI18/MM4_d
+ N_XI45/XI0/NET96_XI45/XI0/XI18/MM4_g N_VSS_XI45/XI0/XI18/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.303e-13
+ PD=5.4e-07 PS=1.45e-06
mXI45/XI0/XI17/MM7 N_XI45/NET273_XI45/XI0/XI17/MM7_d N_NET79_XI45/XI0/XI17/MM7_g
+ N_XI45/XI0/XI17/NET16_XI45/XI0/XI17/MM7_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI17/MM6 N_XI45/XI0/XI17/NET16_XI45/XI0/XI17/MM6_d
+ N_NET95_XI45/XI0/XI17/MM6_g N_XI45/XI0/XI17/NET12_XI45/XI0/XI17/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI17/MM5 N_XI45/XI0/XI17/NET12_XI45/XI0/XI17/MM5_d
+ N_XI45/XI0/NET92_XI45/XI0/XI17/MM5_g N_XI45/XI0/XI17/NET8_XI45/XI0/XI17/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI17/MM4 N_XI45/XI0/XI17/NET8_XI45/XI0/XI17/MM4_d
+ N_XI45/XI0/NET96_XI45/XI0/XI17/MM4_g N_VSS_XI45/XI0/XI17/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.303e-13
+ PD=5.4e-07 PS=1.45e-06
mXI45/XI0/XI16/MM7 N_XI45/NET274_XI45/XI0/XI16/MM7_d N_NET79_XI45/XI0/XI16/MM7_g
+ N_XI45/XI0/XI16/NET16_XI45/XI0/XI16/MM7_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI16/MM6 N_XI45/XI0/XI16/NET16_XI45/XI0/XI16/MM6_d
+ N_XI45/XI0/NET081_XI45/XI0/XI16/MM6_g
+ N_XI45/XI0/XI16/NET12_XI45/XI0/XI16/MM6_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI16/MM5 N_XI45/XI0/XI16/NET12_XI45/XI0/XI16/MM5_d
+ N_NET105_XI45/XI0/XI16/MM5_g N_XI45/XI0/XI16/NET8_XI45/XI0/XI16/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI16/MM4 N_XI45/XI0/XI16/NET8_XI45/XI0/XI16/MM4_d
+ N_XI45/XI0/NET96_XI45/XI0/XI16/MM4_g N_VSS_XI45/XI0/XI16/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.303e-13
+ PD=5.4e-07 PS=1.45e-06
mXI45/XI0/XI15/MM7 N_XI45/NET275_XI45/XI0/XI15/MM7_d N_NET79_XI45/XI0/XI15/MM7_g
+ N_XI45/XI0/XI15/NET16_XI45/XI0/XI15/MM7_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI15/MM6 N_XI45/XI0/XI15/NET16_XI45/XI0/XI15/MM6_d
+ N_NET95_XI45/XI0/XI15/MM6_g N_XI45/XI0/XI15/NET12_XI45/XI0/XI15/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI15/MM5 N_XI45/XI0/XI15/NET12_XI45/XI0/XI15/MM5_d
+ N_NET105_XI45/XI0/XI15/MM5_g N_XI45/XI0/XI15/NET8_XI45/XI0/XI15/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI15/MM4 N_XI45/XI0/XI15/NET8_XI45/XI0/XI15/MM4_d
+ N_XI45/XI0/NET96_XI45/XI0/XI15/MM4_g N_VSS_XI45/XI0/XI15/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.303e-13
+ PD=5.4e-07 PS=1.45e-06
mXI45/XI0/XI14/MM7 N_XI45/NET276_XI45/XI0/XI14/MM7_d N_NET79_XI45/XI0/XI14/MM7_g
+ N_XI45/XI0/XI14/NET16_XI45/XI0/XI14/MM7_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI14/MM6 N_XI45/XI0/XI14/NET16_XI45/XI0/XI14/MM6_d
+ N_XI45/XI0/NET081_XI45/XI0/XI14/MM6_g
+ N_XI45/XI0/XI14/NET12_XI45/XI0/XI14/MM6_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI14/MM5 N_XI45/XI0/XI14/NET12_XI45/XI0/XI14/MM5_d
+ N_XI45/XI0/NET92_XI45/XI0/XI14/MM5_g N_XI45/XI0/XI14/NET8_XI45/XI0/XI14/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI14/MM4 N_XI45/XI0/XI14/NET8_XI45/XI0/XI14/MM4_d
+ N_NET100_XI45/XI0/XI14/MM4_g N_VSS_XI45/XI0/XI14/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.303e-13
+ PD=5.4e-07 PS=1.45e-06
mXI45/XI0/XI13/MM7 N_XI45/NET277_XI45/XI0/XI13/MM7_d N_NET79_XI45/XI0/XI13/MM7_g
+ N_XI45/XI0/XI13/NET16_XI45/XI0/XI13/MM7_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI13/MM6 N_XI45/XI0/XI13/NET16_XI45/XI0/XI13/MM6_d
+ N_NET95_XI45/XI0/XI13/MM6_g N_XI45/XI0/XI13/NET12_XI45/XI0/XI13/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI13/MM5 N_XI45/XI0/XI13/NET12_XI45/XI0/XI13/MM5_d
+ N_XI45/XI0/NET92_XI45/XI0/XI13/MM5_g N_XI45/XI0/XI13/NET8_XI45/XI0/XI13/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI13/MM4 N_XI45/XI0/XI13/NET8_XI45/XI0/XI13/MM4_d
+ N_NET100_XI45/XI0/XI13/MM4_g N_VSS_XI45/XI0/XI13/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.303e-13
+ PD=5.4e-07 PS=1.45e-06
mXI45/XI0/XI12/MM7 N_XI45/NET278_XI45/XI0/XI12/MM7_d N_NET79_XI45/XI0/XI12/MM7_g
+ N_XI45/XI0/XI12/NET16_XI45/XI0/XI12/MM7_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI12/MM6 N_XI45/XI0/XI12/NET16_XI45/XI0/XI12/MM6_d
+ N_XI45/XI0/NET081_XI45/XI0/XI12/MM6_g
+ N_XI45/XI0/XI12/NET12_XI45/XI0/XI12/MM6_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI12/MM5 N_XI45/XI0/XI12/NET12_XI45/XI0/XI12/MM5_d
+ N_NET105_XI45/XI0/XI12/MM5_g N_XI45/XI0/XI12/NET8_XI45/XI0/XI12/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI12/MM4 N_XI45/XI0/XI12/NET8_XI45/XI0/XI12/MM4_d
+ N_NET100_XI45/XI0/XI12/MM4_g N_VSS_XI45/XI0/XI12/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.303e-13
+ PD=5.4e-07 PS=1.45e-06
mXI45/XI0/XI11/MM7 N_XI45/NET266_XI45/XI0/XI11/MM7_d N_NET79_XI45/XI0/XI11/MM7_g
+ N_XI45/XI0/XI11/NET16_XI45/XI0/XI11/MM7_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI11/MM6 N_XI45/XI0/XI11/NET16_XI45/XI0/XI11/MM6_d
+ N_NET95_XI45/XI0/XI11/MM6_g N_XI45/XI0/XI11/NET12_XI45/XI0/XI11/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI11/MM5 N_XI45/XI0/XI11/NET12_XI45/XI0/XI11/MM5_d
+ N_NET105_XI45/XI0/XI11/MM5_g N_XI45/XI0/XI11/NET8_XI45/XI0/XI11/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI11/MM4 N_XI45/XI0/XI11/NET8_XI45/XI0/XI11/MM4_d
+ N_NET100_XI45/XI0/XI11/MM4_g N_VSS_XI45/XI0/XI11/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.303e-13
+ PD=5.4e-07 PS=1.45e-06
mXI45/XI1/XI11/MM4 N_XI45/XI1/XI11/NET8_XI45/XI1/XI11/MM4_d
+ N_NET110_XI45/XI1/XI11/MM4_g N_VSS_XI45/XI1/XI11/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.303e-13
+ PD=5.4e-07 PS=1.45e-06
mXI45/XI1/XI11/MM5 N_XI45/XI1/XI11/NET12_XI45/XI1/XI11/MM5_d
+ N_NET90_XI45/XI1/XI11/MM5_g N_XI45/XI1/XI11/NET8_XI45/XI1/XI11/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI11/MM6 N_XI45/XI1/XI11/NET16_XI45/XI1/XI11/MM6_d
+ N_NET115_XI45/XI1/XI11/MM6_g N_XI45/XI1/XI11/NET12_XI45/XI1/XI11/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI11/MM7 N_XI45/NET252_XI45/XI1/XI11/MM7_d N_NET79_XI45/XI1/XI11/MM7_g
+ N_XI45/XI1/XI11/NET16_XI45/XI1/XI11/MM7_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI12/MM4 N_XI45/XI1/XI12/NET8_XI45/XI1/XI12/MM4_d
+ N_NET110_XI45/XI1/XI12/MM4_g N_VSS_XI45/XI1/XI12/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.303e-13
+ PD=5.4e-07 PS=1.45e-06
mXI45/XI1/XI12/MM5 N_XI45/XI1/XI12/NET12_XI45/XI1/XI12/MM5_d
+ N_NET90_XI45/XI1/XI12/MM5_g N_XI45/XI1/XI12/NET8_XI45/XI1/XI12/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI12/MM6 N_XI45/XI1/XI12/NET16_XI45/XI1/XI12/MM6_d
+ N_XI45/XI1/NET081_XI45/XI1/XI12/MM6_g
+ N_XI45/XI1/XI12/NET12_XI45/XI1/XI12/MM6_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI12/MM7 N_XI45/NET264_XI45/XI1/XI12/MM7_d N_NET79_XI45/XI1/XI12/MM7_g
+ N_XI45/XI1/XI12/NET16_XI45/XI1/XI12/MM7_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI13/MM4 N_XI45/XI1/XI13/NET8_XI45/XI1/XI13/MM4_d
+ N_NET110_XI45/XI1/XI13/MM4_g N_VSS_XI45/XI1/XI13/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.303e-13
+ PD=5.4e-07 PS=1.45e-06
mXI45/XI1/XI13/MM5 N_XI45/XI1/XI13/NET12_XI45/XI1/XI13/MM5_d
+ N_XI45/XI1/NET92_XI45/XI1/XI13/MM5_g N_XI45/XI1/XI13/NET8_XI45/XI1/XI13/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI13/MM6 N_XI45/XI1/XI13/NET16_XI45/XI1/XI13/MM6_d
+ N_NET115_XI45/XI1/XI13/MM6_g N_XI45/XI1/XI13/NET12_XI45/XI1/XI13/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI13/MM7 N_XI45/NET263_XI45/XI1/XI13/MM7_d N_NET79_XI45/XI1/XI13/MM7_g
+ N_XI45/XI1/XI13/NET16_XI45/XI1/XI13/MM7_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI14/MM4 N_XI45/XI1/XI14/NET8_XI45/XI1/XI14/MM4_d
+ N_NET110_XI45/XI1/XI14/MM4_g N_VSS_XI45/XI1/XI14/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.303e-13
+ PD=5.4e-07 PS=1.45e-06
mXI45/XI1/XI14/MM5 N_XI45/XI1/XI14/NET12_XI45/XI1/XI14/MM5_d
+ N_XI45/XI1/NET92_XI45/XI1/XI14/MM5_g N_XI45/XI1/XI14/NET8_XI45/XI1/XI14/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI14/MM6 N_XI45/XI1/XI14/NET16_XI45/XI1/XI14/MM6_d
+ N_XI45/XI1/NET081_XI45/XI1/XI14/MM6_g
+ N_XI45/XI1/XI14/NET12_XI45/XI1/XI14/MM6_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI14/MM7 N_XI45/NET262_XI45/XI1/XI14/MM7_d N_NET79_XI45/XI1/XI14/MM7_g
+ N_XI45/XI1/XI14/NET16_XI45/XI1/XI14/MM7_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI15/MM4 N_XI45/XI1/XI15/NET8_XI45/XI1/XI15/MM4_d
+ N_XI45/XI1/NET96_XI45/XI1/XI15/MM4_g N_VSS_XI45/XI1/XI15/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.303e-13
+ PD=5.4e-07 PS=1.45e-06
mXI45/XI1/XI15/MM5 N_XI45/XI1/XI15/NET12_XI45/XI1/XI15/MM5_d
+ N_NET90_XI45/XI1/XI15/MM5_g N_XI45/XI1/XI15/NET8_XI45/XI1/XI15/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI15/MM6 N_XI45/XI1/XI15/NET16_XI45/XI1/XI15/MM6_d
+ N_NET115_XI45/XI1/XI15/MM6_g N_XI45/XI1/XI15/NET12_XI45/XI1/XI15/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI15/MM7 N_XI45/NET261_XI45/XI1/XI15/MM7_d N_NET79_XI45/XI1/XI15/MM7_g
+ N_XI45/XI1/XI15/NET16_XI45/XI1/XI15/MM7_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI16/MM4 N_XI45/XI1/XI16/NET8_XI45/XI1/XI16/MM4_d
+ N_XI45/XI1/NET96_XI45/XI1/XI16/MM4_g N_VSS_XI45/XI1/XI16/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.303e-13
+ PD=5.4e-07 PS=1.45e-06
mXI45/XI1/XI16/MM5 N_XI45/XI1/XI16/NET12_XI45/XI1/XI16/MM5_d
+ N_NET90_XI45/XI1/XI16/MM5_g N_XI45/XI1/XI16/NET8_XI45/XI1/XI16/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI16/MM6 N_XI45/XI1/XI16/NET16_XI45/XI1/XI16/MM6_d
+ N_XI45/XI1/NET081_XI45/XI1/XI16/MM6_g
+ N_XI45/XI1/XI16/NET12_XI45/XI1/XI16/MM6_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI16/MM7 N_XI45/NET260_XI45/XI1/XI16/MM7_d N_NET79_XI45/XI1/XI16/MM7_g
+ N_XI45/XI1/XI16/NET16_XI45/XI1/XI16/MM7_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI17/MM4 N_XI45/XI1/XI17/NET8_XI45/XI1/XI17/MM4_d
+ N_XI45/XI1/NET96_XI45/XI1/XI17/MM4_g N_VSS_XI45/XI1/XI17/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.303e-13
+ PD=5.4e-07 PS=1.45e-06
mXI45/XI1/XI17/MM5 N_XI45/XI1/XI17/NET12_XI45/XI1/XI17/MM5_d
+ N_XI45/XI1/NET92_XI45/XI1/XI17/MM5_g N_XI45/XI1/XI17/NET8_XI45/XI1/XI17/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI17/MM6 N_XI45/XI1/XI17/NET16_XI45/XI1/XI17/MM6_d
+ N_NET115_XI45/XI1/XI17/MM6_g N_XI45/XI1/XI17/NET12_XI45/XI1/XI17/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI17/MM7 N_XI45/NET259_XI45/XI1/XI17/MM7_d N_NET79_XI45/XI1/XI17/MM7_g
+ N_XI45/XI1/XI17/NET16_XI45/XI1/XI17/MM7_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI18/MM4 N_XI45/XI1/XI18/NET8_XI45/XI1/XI18/MM4_d
+ N_XI45/XI1/NET96_XI45/XI1/XI18/MM4_g N_VSS_XI45/XI1/XI18/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.303e-13
+ PD=5.4e-07 PS=1.45e-06
mXI45/XI1/XI18/MM5 N_XI45/XI1/XI18/NET12_XI45/XI1/XI18/MM5_d
+ N_XI45/XI1/NET92_XI45/XI1/XI18/MM5_g N_XI45/XI1/XI18/NET8_XI45/XI1/XI18/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI18/MM6 N_XI45/XI1/XI18/NET16_XI45/XI1/XI18/MM6_d
+ N_XI45/XI1/NET081_XI45/XI1/XI18/MM6_g
+ N_XI45/XI1/XI18/NET12_XI45/XI1/XI18/MM6_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI18/MM7 N_XI45/NET258_XI45/XI1/XI18/MM7_d N_NET79_XI45/XI1/XI18/MM7_g
+ N_XI45/XI1/XI18/NET16_XI45/XI1/XI18/MM7_s N_VSS_XI45/XI0/XI8/MM0_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI47/MM3 N_NET0215_XI47/MM3_d N_NET0265_XI47/MM3_g N_DOUT<0>_XI47/MM3_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=7.5e-07 AD=3.675e-13 AS=1.92e-13
+ PD=1.73e-06 PS=8.58e-07
mXI47/MM0 N_NET0214_XI47/MM0_d N_NET0265_XI47/MM0_g N_NET0183_XI47/MM0_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=7.5e-07 AD=3.675e-13 AS=1.92e-13
+ PD=1.73e-06 PS=8.58e-07
mXI47/MM1 N_DOUT<0>_XI47/MM1_d N_NET0183_XI47/MM1_g N_VSS_XI47/MM1_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.28e-13 AS=1.8e-13
+ PD=5.72e-07 PS=7.2e-07
mXI47/MM2 N_NET0183_XI47/MM2_d N_DOUT<0>_XI47/MM2_g N_VSS_XI47/MM2_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.28e-13 AS=1.8e-13
+ PD=5.72e-07 PS=7.2e-07
mXI19/MM7 N_XI19/NET0139_XI19/MM7_d N_XI19/NET41_XI19/MM7_g N_VSS_XI19/MM7_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI19/MM4 N_XI19/NET41_XI19/MM4_d N_CLK_XI19/MM4_g N_VSS_XI19/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI19/MM2 N_NET81_XI19/MM2_d N_XI19/NET49_XI19/MM2_g N_VSS_XI19/MM2_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI19/MM1 N_XI19/NET49_XI19/MM1_d N_CLK_XI19/MM1_g N_VSS_XI19/MM1_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI11/MM7 N_XI11/NET13_XI11/MM7_d N_A<8>_XI11/MM7_g N_VSS_XI11/MM7_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI11/MM8 N_XI11/NET9_XI11/MM8_d N_CLK_XI11/MM8_g N_VSS_XI11/MM8_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI11/MM5 N_XI11/NET21_XI11/MM5_d N_XI11/NET13_XI11/MM5_g N_XI11/NET9_XI11/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI11/MM9 N_XI11/NET5_XI11/MM9_d N_XI11/NET21_XI11/MM9_g N_VSS_XI11/MM9_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI11/MM6 N_XI11/NET15_XI11/MM6_d N_CLK_XI11/MM6_g N_XI11/NET5_XI11/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI11/MM10 N_NET120_XI11/MM10_d N_XI11/NET15_XI11/MM10_g N_VSS_XI11/MM10_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI12/MM7 N_XI12/NET13_XI12/MM7_d N_A<5>_XI12/MM7_g N_VSS_XI12/MM7_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI12/MM8 N_XI12/NET9_XI12/MM8_d N_CLK_XI12/MM8_g N_VSS_XI12/MM8_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI12/MM5 N_XI12/NET21_XI12/MM5_d N_XI12/NET13_XI12/MM5_g N_XI12/NET9_XI12/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI12/MM9 N_XI12/NET5_XI12/MM9_d N_XI12/NET21_XI12/MM9_g N_VSS_XI12/MM9_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI12/MM6 N_XI12/NET15_XI12/MM6_d N_CLK_XI12/MM6_g N_XI12/NET5_XI12/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI12/MM10 N_NET115_XI12/MM10_d N_XI12/NET15_XI12/MM10_g N_VSS_XI12/MM10_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI17/MM7 N_XI17/NET13_XI17/MM7_d N_A<4>_XI17/MM7_g N_VSS_XI17/MM7_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI17/MM8 N_XI17/NET9_XI17/MM8_d N_CLK_XI17/MM8_g N_VSS_XI17/MM8_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI17/MM5 N_XI17/NET21_XI17/MM5_d N_XI17/NET13_XI17/MM5_g N_XI17/NET9_XI17/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI17/MM9 N_XI17/NET5_XI17/MM9_d N_XI17/NET21_XI17/MM9_g N_VSS_XI17/MM9_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI17/MM6 N_XI17/NET15_XI17/MM6_d N_CLK_XI17/MM6_g N_XI17/NET5_XI17/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI17/MM10 N_NET90_XI17/MM10_d N_XI17/NET15_XI17/MM10_g N_VSS_XI17/MM10_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI13/MM7 N_XI13/NET13_XI13/MM7_d N_A<3>_XI13/MM7_g N_VSS_XI13/MM7_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI13/MM8 N_XI13/NET9_XI13/MM8_d N_CLK_XI13/MM8_g N_VSS_XI13/MM8_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI13/MM5 N_XI13/NET21_XI13/MM5_d N_XI13/NET13_XI13/MM5_g N_XI13/NET9_XI13/MM5_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI13/MM9 N_XI13/NET5_XI13/MM9_d N_XI13/NET21_XI13/MM9_g N_VSS_XI13/MM9_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=5.875e-14 AS=2.303e-13
+ PD=2.5e-07 PS=1.45e-06
mXI13/MM6 N_XI13/NET15_XI13/MM6_d N_CLK_XI13/MM6_g N_XI13/NET5_XI13/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=5.875e-14
+ PD=1.45e-06 PS=2.5e-07
mXI13/MM10 N_NET110_XI13/MM10_d N_XI13/NET15_XI13/MM10_g N_VSS_XI13/MM10_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI19/MM18 N_XI19/NET37_XI19/MM18_d N_XI19/NET0139_XI19/MM18_g N_VSS_XI19/MM18_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI19/XI0/MM3 N_XI19/XI0/NET5_XI19/XI0/MM3_d N_XI19/NET37_XI19/XI0/MM3_g
+ N_VSS_XI19/XI0/MM3_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06
mXI19/XI0/MM2 N_NET79_XI19/XI0/MM2_d N_NET81_XI19/XI0/MM2_g
+ N_XI19/XI0/NET5_XI19/XI0/MM2_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.6685e-13 PD=1.45e-06 PS=7.1e-07
mXI19/MM22 N_XI19/NET082_XI19/MM22_d N_NET81_XI19/MM22_g N_VSS_XI19/MM22_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI19/MM21 N_XI19/NET086_XI19/MM21_d N_XI19/NET082_XI19/MM21_g N_VSS_XI19/MM21_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=3e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI19/MM25 N_NET0265_XI19/MM25_d N_XI19/NET0100_XI19/MM25_g N_VSS_XI19/MM25_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI19/MM28 N_XI19/NET0100_XI19/MM28_d N_NET82_XI19/MM28_g N_VSS_XI19/MM28_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.773e-13
+ PD=1.45e-06 PS=1.65e-06
mXI19/MM16 N_NET82_XI19/MM16_d N_XI19/NET9_XI19/MM16_g N_VSS_XI19/MM16_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI19/XI1/MM2 N_XI19/NET9_XI19/XI1/MM2_d N_XI19/NET086_XI19/XI1/MM2_g
+ N_XI19/XI1/NET5_XI19/XI1/MM2_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.6685e-13 PD=1.45e-06 PS=7.1e-07
mXI19/XI1/MM3 N_XI19/XI1/NET5_XI19/XI1/MM3_d N_XI19/NET086_XI19/XI1/MM3_g
+ N_VSS_XI19/XI1/MM3_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06
mXI49/MM0 N_NET0208_XI49/MM0_d N_NET0207_XI49/MM0_g N_VSS_XI49/MM0_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI48/MM0 N_NET0207_XI48/MM0_d N_NET141_XI48/MM0_g N_VSS_XI48/MM0_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI8/MM1 N_NET141_XI8/MM1_d N_NET0174_XI8/MM1_g N_XI8/NET40_XI8/MM1_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=1e-06 AD=5e-13 AS=1.5e-13 PD=2e-06
+ PS=3e-07
mXI8/MM0 N_XI8/NET40_XI8/MM0_d N_VREF_XI8/MM0_g N_XI8/NET43_XI8/MM0_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=1e-06 AD=1.5e-13 AS=2.7e-13 PD=3e-07
+ PS=5.4e-07
mXI8/MM4 N_XI8/NET43_XI8/MM4_d N_NET82_XI8/MM4_g N_VSS_XI8/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=1e-06 AD=2.7e-13 AS=2.55e-13
+ PD=5.4e-07 PS=5.1e-07
mXI8/MM4@2 N_XI8/NET43_XI8/MM4@2_d N_NET82_XI8/MM4@2_g N_VSS_XI8/MM4@2_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=1e-06 AD=2.7e-13 AS=2.55e-13
+ PD=5.4e-07 PS=5.1e-07
mXI8/MM3 N_XI8/NET28_XI8/MM3_d N_NET139_XI8/MM3_g N_XI8/NET43_XI8/MM3_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=1e-06 AD=1.725e-13 AS=2.7e-13
+ PD=3.45e-07 PS=5.4e-07
mXI8/MM2 N_NET0174_XI8/MM2_d N_NET141_XI8/MM2_g N_XI8/NET28_XI8/MM2_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=1.725e-13
+ PD=1.98e-06 PS=3.45e-07
mXI45/XI58/MM1 N_NET10_XI45/XI58/MM1_d N_XI45/NET272_XI45/XI58/MM1_g
+ N_VSS_XI45/XI58/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI59/MM1 N_NET11_XI45/XI59/MM1_d N_XI45/NET272_XI45/XI59/MM1_g
+ N_VSS_XI45/XI59/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI60/MM1 N_NET12_XI45/XI60/MM1_d N_XI45/NET272_XI45/XI60/MM1_g
+ N_VSS_XI45/XI60/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI61/MM1 N_NET13_XI45/XI61/MM1_d N_XI45/NET272_XI45/XI61/MM1_g
+ N_VSS_XI45/XI61/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI62/MM1 N_NET14_XI45/XI62/MM1_d N_XI45/NET272_XI45/XI62/MM1_g
+ N_VSS_XI45/XI62/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI63/MM1 N_NET15_XI45/XI63/MM1_d N_XI45/NET272_XI45/XI63/MM1_g
+ N_VSS_XI45/XI63/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI64/MM1 N_NET16_XI45/XI64/MM1_d N_XI45/NET272_XI45/XI64/MM1_g
+ N_VSS_XI45/XI64/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI65/MM1 N_NET17_XI45/XI65/MM1_d N_XI45/NET272_XI45/XI65/MM1_g
+ N_VSS_XI45/XI65/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI57/MM1 N_NET18_XI45/XI57/MM1_d N_XI45/NET273_XI45/XI57/MM1_g
+ N_VSS_XI45/XI57/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI56/MM1 N_NET19_XI45/XI56/MM1_d N_XI45/NET273_XI45/XI56/MM1_g
+ N_VSS_XI45/XI56/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI55/MM1 N_NET20_XI45/XI55/MM1_d N_XI45/NET273_XI45/XI55/MM1_g
+ N_VSS_XI45/XI55/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI54/MM1 N_NET21_XI45/XI54/MM1_d N_XI45/NET273_XI45/XI54/MM1_g
+ N_VSS_XI45/XI54/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI53/MM1 N_NET22_XI45/XI53/MM1_d N_XI45/NET273_XI45/XI53/MM1_g
+ N_VSS_XI45/XI53/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI52/MM1 N_NET23_XI45/XI52/MM1_d N_XI45/NET273_XI45/XI52/MM1_g
+ N_VSS_XI45/XI52/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI51/MM1 N_NET24_XI45/XI51/MM1_d N_XI45/NET273_XI45/XI51/MM1_g
+ N_VSS_XI45/XI51/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI50/MM1 N_NET25_XI45/XI50/MM1_d N_XI45/NET273_XI45/XI50/MM1_g
+ N_VSS_XI45/XI50/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI42/MM1 N_NET26_XI45/XI42/MM1_d N_XI45/NET274_XI45/XI42/MM1_g
+ N_VSS_XI45/XI42/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI43/MM1 N_NET27_XI45/XI43/MM1_d N_XI45/NET274_XI45/XI43/MM1_g
+ N_VSS_XI45/XI43/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI44/MM1 N_NET28_XI45/XI44/MM1_d N_XI45/NET274_XI45/XI44/MM1_g
+ N_VSS_XI45/XI44/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI45/MM1 N_NET29_XI45/XI45/MM1_d N_XI45/NET274_XI45/XI45/MM1_g
+ N_VSS_XI45/XI45/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI46/MM1 N_NET30_XI45/XI46/MM1_d N_XI45/NET274_XI45/XI46/MM1_g
+ N_VSS_XI45/XI46/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI47/MM1 N_NET31_XI45/XI47/MM1_d N_XI45/NET274_XI45/XI47/MM1_g
+ N_VSS_XI45/XI47/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI48/MM1 N_NET32_XI45/XI48/MM1_d N_XI45/NET274_XI45/XI48/MM1_g
+ N_VSS_XI45/XI48/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI49/MM1 N_NET33_XI45/XI49/MM1_d N_XI45/NET274_XI45/XI49/MM1_g
+ N_VSS_XI45/XI49/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI41/MM1 N_NET34_XI45/XI41/MM1_d N_XI45/NET275_XI45/XI41/MM1_g
+ N_VSS_XI45/XI41/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI40/MM1 N_NET35_XI45/XI40/MM1_d N_XI45/NET275_XI45/XI40/MM1_g
+ N_VSS_XI45/XI40/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI39/MM1 N_NET36_XI45/XI39/MM1_d N_XI45/NET275_XI45/XI39/MM1_g
+ N_VSS_XI45/XI39/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI38/MM1 N_NET37_XI45/XI38/MM1_d N_XI45/NET275_XI45/XI38/MM1_g
+ N_VSS_XI45/XI38/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI37/MM1 N_NET38_XI45/XI37/MM1_d N_XI45/NET275_XI45/XI37/MM1_g
+ N_VSS_XI45/XI37/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI36/MM1 N_NET39_XI45/XI36/MM1_d N_XI45/NET275_XI45/XI36/MM1_g
+ N_VSS_XI45/XI36/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI35/MM1 N_NET40_XI45/XI35/MM1_d N_XI45/NET275_XI45/XI35/MM1_g
+ N_VSS_XI45/XI35/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI34/MM1 N_NET41_XI45/XI34/MM1_d N_XI45/NET275_XI45/XI34/MM1_g
+ N_VSS_XI45/XI34/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI26/MM1 N_NET42_XI45/XI26/MM1_d N_XI45/NET276_XI45/XI26/MM1_g
+ N_VSS_XI45/XI26/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI27/MM1 N_NET43_XI45/XI27/MM1_d N_XI45/NET276_XI45/XI27/MM1_g
+ N_VSS_XI45/XI27/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI28/MM1 N_NET44_XI45/XI28/MM1_d N_XI45/NET276_XI45/XI28/MM1_g
+ N_VSS_XI45/XI28/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI29/MM1 N_NET45_XI45/XI29/MM1_d N_XI45/NET276_XI45/XI29/MM1_g
+ N_VSS_XI45/XI29/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI30/MM1 N_NET46_XI45/XI30/MM1_d N_XI45/NET276_XI45/XI30/MM1_g
+ N_VSS_XI45/XI30/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI31/MM1 N_NET47_XI45/XI31/MM1_d N_XI45/NET276_XI45/XI31/MM1_g
+ N_VSS_XI45/XI31/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI32/MM1 N_NET48_XI45/XI32/MM1_d N_XI45/NET276_XI45/XI32/MM1_g
+ N_VSS_XI45/XI32/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI33/MM1 N_NET49_XI45/XI33/MM1_d N_XI45/NET276_XI45/XI33/MM1_g
+ N_VSS_XI45/XI33/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI25/MM1 N_NET50_XI45/XI25/MM1_d N_XI45/NET277_XI45/XI25/MM1_g
+ N_VSS_XI45/XI25/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI24/MM1 N_NET51_XI45/XI24/MM1_d N_XI45/NET277_XI45/XI24/MM1_g
+ N_VSS_XI45/XI24/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI23/MM1 N_NET52_XI45/XI23/MM1_d N_XI45/NET277_XI45/XI23/MM1_g
+ N_VSS_XI45/XI23/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI22/MM1 N_NET53_XI45/XI22/MM1_d N_XI45/NET277_XI45/XI22/MM1_g
+ N_VSS_XI45/XI22/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI21/MM1 N_NET54_XI45/XI21/MM1_d N_XI45/NET277_XI45/XI21/MM1_g
+ N_VSS_XI45/XI21/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI20/MM1 N_NET55_XI45/XI20/MM1_d N_XI45/NET277_XI45/XI20/MM1_g
+ N_VSS_XI45/XI20/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI19/MM1 N_NET56_XI45/XI19/MM1_d N_XI45/NET277_XI45/XI19/MM1_g
+ N_VSS_XI45/XI19/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI18/MM1 N_NET57_XI45/XI18/MM1_d N_XI45/NET277_XI45/XI18/MM1_g
+ N_VSS_XI45/XI18/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI10/MM1 N_NET58_XI45/XI10/MM1_d N_XI45/NET278_XI45/XI10/MM1_g
+ N_VSS_XI45/XI10/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI11/MM1 N_NET59_XI45/XI11/MM1_d N_XI45/NET278_XI45/XI11/MM1_g
+ N_VSS_XI45/XI11/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI12/MM1 N_NET60_XI45/XI12/MM1_d N_XI45/NET278_XI45/XI12/MM1_g
+ N_VSS_XI45/XI12/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI13/MM1 N_NET61_XI45/XI13/MM1_d N_XI45/NET278_XI45/XI13/MM1_g
+ N_VSS_XI45/XI13/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI14/MM1 N_NET62_XI45/XI14/MM1_d N_XI45/NET278_XI45/XI14/MM1_g
+ N_VSS_XI45/XI14/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI15/MM1 N_NET63_XI45/XI15/MM1_d N_XI45/NET278_XI45/XI15/MM1_g
+ N_VSS_XI45/XI15/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI16/MM1 N_NET64_XI45/XI16/MM1_d N_XI45/NET278_XI45/XI16/MM1_g
+ N_VSS_XI45/XI16/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI17/MM1 N_NET65_XI45/XI17/MM1_d N_XI45/NET278_XI45/XI17/MM1_g
+ N_VSS_XI45/XI17/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI9/MM1 N_NET66_XI45/XI9/MM1_d N_XI45/NET266_XI45/XI9/MM1_g
+ N_VSS_XI45/XI9/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI8/MM1 N_NET67_XI45/XI8/MM1_d N_XI45/NET266_XI45/XI8/MM1_g
+ N_VSS_XI45/XI8/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI7/MM1 N_NET68_XI45/XI7/MM1_d N_XI45/NET266_XI45/XI7/MM1_g
+ N_VSS_XI45/XI7/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI6/MM1 N_NET69_XI45/XI6/MM1_d N_XI45/NET266_XI45/XI6/MM1_g
+ N_VSS_XI45/XI6/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI5/MM1 N_NET70_XI45/XI5/MM1_d N_XI45/NET266_XI45/XI5/MM1_g
+ N_VSS_XI45/XI5/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI4/MM1 N_NET71_XI45/XI4/MM1_d N_XI45/NET266_XI45/XI4/MM1_g
+ N_VSS_XI45/XI4/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI3/MM1 N_NET72_XI45/XI3/MM1_d N_XI45/NET266_XI45/XI3/MM1_g
+ N_VSS_XI45/XI3/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI2/MM1 N_NET8_XI45/XI2/MM1_d N_XI45/NET266_XI45/XI2/MM1_g
+ N_VSS_XI45/XI2/MM1_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI7/MM4 N_XI7/NET48_XI7/MM4_d N_NET120_XI7/MM4_g N_VSS_XI7/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI45/XI58/MM0 N_NET10_XI45/XI58/MM0_d N_XI45/NET258_XI45/XI58/MM0_g
+ N_VSS_XI45/XI58/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI59/MM0 N_NET11_XI45/XI59/MM0_d N_XI45/NET259_XI45/XI59/MM0_g
+ N_VSS_XI45/XI59/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI60/MM0 N_NET12_XI45/XI60/MM0_d N_XI45/NET260_XI45/XI60/MM0_g
+ N_VSS_XI45/XI60/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI61/MM0 N_NET13_XI45/XI61/MM0_d N_XI45/NET261_XI45/XI61/MM0_g
+ N_VSS_XI45/XI61/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI62/MM0 N_NET14_XI45/XI62/MM0_d N_XI45/NET262_XI45/XI62/MM0_g
+ N_VSS_XI45/XI62/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI63/MM0 N_NET15_XI45/XI63/MM0_d N_XI45/NET263_XI45/XI63/MM0_g
+ N_VSS_XI45/XI63/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI64/MM0 N_NET16_XI45/XI64/MM0_d N_XI45/NET264_XI45/XI64/MM0_g
+ N_VSS_XI45/XI64/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI65/MM0 N_NET17_XI45/XI65/MM0_d N_XI45/NET252_XI45/XI65/MM0_g
+ N_VSS_XI45/XI65/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI57/MM0 N_NET18_XI45/XI57/MM0_d N_XI45/NET258_XI45/XI57/MM0_g
+ N_VSS_XI45/XI57/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI56/MM0 N_NET19_XI45/XI56/MM0_d N_XI45/NET259_XI45/XI56/MM0_g
+ N_VSS_XI45/XI56/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI55/MM0 N_NET20_XI45/XI55/MM0_d N_XI45/NET260_XI45/XI55/MM0_g
+ N_VSS_XI45/XI55/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI54/MM0 N_NET21_XI45/XI54/MM0_d N_XI45/NET261_XI45/XI54/MM0_g
+ N_VSS_XI45/XI54/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI53/MM0 N_NET22_XI45/XI53/MM0_d N_XI45/NET262_XI45/XI53/MM0_g
+ N_VSS_XI45/XI53/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI52/MM0 N_NET23_XI45/XI52/MM0_d N_XI45/NET263_XI45/XI52/MM0_g
+ N_VSS_XI45/XI52/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI51/MM0 N_NET24_XI45/XI51/MM0_d N_XI45/NET264_XI45/XI51/MM0_g
+ N_VSS_XI45/XI51/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI50/MM0 N_NET25_XI45/XI50/MM0_d N_XI45/NET252_XI45/XI50/MM0_g
+ N_VSS_XI45/XI50/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI42/MM0 N_NET26_XI45/XI42/MM0_d N_XI45/NET258_XI45/XI42/MM0_g
+ N_VSS_XI45/XI42/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI43/MM0 N_NET27_XI45/XI43/MM0_d N_XI45/NET259_XI45/XI43/MM0_g
+ N_VSS_XI45/XI43/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI44/MM0 N_NET28_XI45/XI44/MM0_d N_XI45/NET260_XI45/XI44/MM0_g
+ N_VSS_XI45/XI44/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI45/MM0 N_NET29_XI45/XI45/MM0_d N_XI45/NET261_XI45/XI45/MM0_g
+ N_VSS_XI45/XI45/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI46/MM0 N_NET30_XI45/XI46/MM0_d N_XI45/NET262_XI45/XI46/MM0_g
+ N_VSS_XI45/XI46/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI47/MM0 N_NET31_XI45/XI47/MM0_d N_XI45/NET263_XI45/XI47/MM0_g
+ N_VSS_XI45/XI47/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI48/MM0 N_NET32_XI45/XI48/MM0_d N_XI45/NET264_XI45/XI48/MM0_g
+ N_VSS_XI45/XI48/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI49/MM0 N_NET33_XI45/XI49/MM0_d N_XI45/NET252_XI45/XI49/MM0_g
+ N_VSS_XI45/XI49/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI41/MM0 N_NET34_XI45/XI41/MM0_d N_XI45/NET258_XI45/XI41/MM0_g
+ N_VSS_XI45/XI41/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI40/MM0 N_NET35_XI45/XI40/MM0_d N_XI45/NET259_XI45/XI40/MM0_g
+ N_VSS_XI45/XI40/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI39/MM0 N_NET36_XI45/XI39/MM0_d N_XI45/NET260_XI45/XI39/MM0_g
+ N_VSS_XI45/XI39/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI38/MM0 N_NET37_XI45/XI38/MM0_d N_XI45/NET261_XI45/XI38/MM0_g
+ N_VSS_XI45/XI38/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI37/MM0 N_NET38_XI45/XI37/MM0_d N_XI45/NET262_XI45/XI37/MM0_g
+ N_VSS_XI45/XI37/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI36/MM0 N_NET39_XI45/XI36/MM0_d N_XI45/NET263_XI45/XI36/MM0_g
+ N_VSS_XI45/XI36/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI35/MM0 N_NET40_XI45/XI35/MM0_d N_XI45/NET264_XI45/XI35/MM0_g
+ N_VSS_XI45/XI35/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI34/MM0 N_NET41_XI45/XI34/MM0_d N_XI45/NET252_XI45/XI34/MM0_g
+ N_VSS_XI45/XI34/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI26/MM0 N_NET42_XI45/XI26/MM0_d N_XI45/NET258_XI45/XI26/MM0_g
+ N_VSS_XI45/XI26/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI27/MM0 N_NET43_XI45/XI27/MM0_d N_XI45/NET259_XI45/XI27/MM0_g
+ N_VSS_XI45/XI27/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI28/MM0 N_NET44_XI45/XI28/MM0_d N_XI45/NET260_XI45/XI28/MM0_g
+ N_VSS_XI45/XI28/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI29/MM0 N_NET45_XI45/XI29/MM0_d N_XI45/NET261_XI45/XI29/MM0_g
+ N_VSS_XI45/XI29/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI30/MM0 N_NET46_XI45/XI30/MM0_d N_XI45/NET262_XI45/XI30/MM0_g
+ N_VSS_XI45/XI30/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI31/MM0 N_NET47_XI45/XI31/MM0_d N_XI45/NET263_XI45/XI31/MM0_g
+ N_VSS_XI45/XI31/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI32/MM0 N_NET48_XI45/XI32/MM0_d N_XI45/NET264_XI45/XI32/MM0_g
+ N_VSS_XI45/XI32/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI33/MM0 N_NET49_XI45/XI33/MM0_d N_XI45/NET252_XI45/XI33/MM0_g
+ N_VSS_XI45/XI33/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI25/MM0 N_NET50_XI45/XI25/MM0_d N_XI45/NET258_XI45/XI25/MM0_g
+ N_VSS_XI45/XI25/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI24/MM0 N_NET51_XI45/XI24/MM0_d N_XI45/NET259_XI45/XI24/MM0_g
+ N_VSS_XI45/XI24/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI23/MM0 N_NET52_XI45/XI23/MM0_d N_XI45/NET260_XI45/XI23/MM0_g
+ N_VSS_XI45/XI23/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI22/MM0 N_NET53_XI45/XI22/MM0_d N_XI45/NET261_XI45/XI22/MM0_g
+ N_VSS_XI45/XI22/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI21/MM0 N_NET54_XI45/XI21/MM0_d N_XI45/NET262_XI45/XI21/MM0_g
+ N_VSS_XI45/XI21/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI20/MM0 N_NET55_XI45/XI20/MM0_d N_XI45/NET263_XI45/XI20/MM0_g
+ N_VSS_XI45/XI20/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI19/MM0 N_NET56_XI45/XI19/MM0_d N_XI45/NET264_XI45/XI19/MM0_g
+ N_VSS_XI45/XI19/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI18/MM0 N_NET57_XI45/XI18/MM0_d N_XI45/NET252_XI45/XI18/MM0_g
+ N_VSS_XI45/XI18/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI10/MM0 N_NET58_XI45/XI10/MM0_d N_XI45/NET258_XI45/XI10/MM0_g
+ N_VSS_XI45/XI10/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI11/MM0 N_NET59_XI45/XI11/MM0_d N_XI45/NET259_XI45/XI11/MM0_g
+ N_VSS_XI45/XI11/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI12/MM0 N_NET60_XI45/XI12/MM0_d N_XI45/NET260_XI45/XI12/MM0_g
+ N_VSS_XI45/XI12/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI13/MM0 N_NET61_XI45/XI13/MM0_d N_XI45/NET261_XI45/XI13/MM0_g
+ N_VSS_XI45/XI13/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI14/MM0 N_NET62_XI45/XI14/MM0_d N_XI45/NET262_XI45/XI14/MM0_g
+ N_VSS_XI45/XI14/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI15/MM0 N_NET63_XI45/XI15/MM0_d N_XI45/NET263_XI45/XI15/MM0_g
+ N_VSS_XI45/XI15/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI16/MM0 N_NET64_XI45/XI16/MM0_d N_XI45/NET264_XI45/XI16/MM0_g
+ N_VSS_XI45/XI16/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI17/MM0 N_NET65_XI45/XI17/MM0_d N_XI45/NET252_XI45/XI17/MM0_g
+ N_VSS_XI45/XI17/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI9/MM0 N_NET66_XI45/XI9/MM0_d N_XI45/NET258_XI45/XI9/MM0_g
+ N_VSS_XI45/XI9/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI8/MM0 N_NET67_XI45/XI8/MM0_d N_XI45/NET259_XI45/XI8/MM0_g
+ N_VSS_XI45/XI8/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI7/MM0 N_NET68_XI45/XI7/MM0_d N_XI45/NET260_XI45/XI7/MM0_g
+ N_VSS_XI45/XI7/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI6/MM0 N_NET69_XI45/XI6/MM0_d N_XI45/NET261_XI45/XI6/MM0_g
+ N_VSS_XI45/XI6/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI5/MM0 N_NET70_XI45/XI5/MM0_d N_XI45/NET262_XI45/XI5/MM0_g
+ N_VSS_XI45/XI5/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI4/MM0 N_NET71_XI45/XI4/MM0_d N_XI45/NET263_XI45/XI4/MM0_g
+ N_VSS_XI45/XI4/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI3/MM0 N_NET72_XI45/XI3/MM0_d N_XI45/NET264_XI45/XI3/MM0_g
+ N_VSS_XI45/XI3/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI45/XI2/MM0 N_NET8_XI45/XI2/MM0_d N_XI45/NET252_XI45/XI2/MM0_g
+ N_VSS_XI45/XI2/MM0_s N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI7/MM6 N_XI7/NET68_XI7/MM6_d N_NET125_XI7/MM6_g N_VSS_XI7/MM6_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI7/MM9 N_XI7/NET76_XI7/MM9_d N_NET85_XI7/MM9_g N_VSS_XI7/MM9_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI7/MM1 N_NET147_XI7/MM1_d N_NET120_XI7/MM1_g N_XI7/NET141_XI7/MM1_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI5/MM1040 N_NET147_XI5/MM1040_d N_NET10_XI5/MM1040_g N_VSS_XI5/MM1040_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1332 XI5/NET02326 N_NET11_XI5/MM1332_g N_VSS_XI5/MM1332_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1039 N_NET147_XI5/MM1039_d N_NET12_XI5/MM1039_g N_VSS_XI5/MM1039_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1321 XI5/NET02370 N_NET13_XI5/MM1321_g N_VSS_XI5/MM1321_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1008 N_NET147_XI5/MM1008_d N_NET14_XI5/MM1008_g N_VSS_XI5/MM1008_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1313 XI5/NET02402 N_NET15_XI5/MM1313_g N_VSS_XI5/MM1313_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1007 N_NET147_XI5/MM1007_d N_NET16_XI5/MM1007_g N_VSS_XI5/MM1007_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1305 XI5/NET02434 N_NET17_XI5/MM1305_g N_VSS_XI5/MM1305_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM976 N_NET147_XI5/MM976_d N_NET18_XI5/MM976_g N_VSS_XI5/MM976_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1297 XI5/NET02466 N_NET19_XI5/MM1297_g N_VSS_XI5/MM1297_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM975 N_NET147_XI5/MM975_d N_NET20_XI5/MM975_g N_VSS_XI5/MM975_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1289 XI5/NET04286 N_NET21_XI5/MM1289_g N_VSS_XI5/MM1289_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM944 N_NET147_XI5/MM944_d N_NET22_XI5/MM944_g N_VSS_XI5/MM944_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1281 XI5/NET04318 N_NET23_XI5/MM1281_g N_VSS_XI5/MM1281_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM943 N_NET147_XI5/MM943_d N_NET24_XI5/MM943_g N_VSS_XI5/MM943_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1273 XI5/NET03466 N_NET25_XI5/MM1273_g N_VSS_XI5/MM1273_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM912 N_NET147_XI5/MM912_d N_NET26_XI5/MM912_g N_VSS_XI5/MM912_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1272 XI5/NET05406 N_NET27_XI5/MM1272_g N_VSS_XI5/MM1272_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM911 N_NET147_XI5/MM911_d N_NET28_XI5/MM911_g N_VSS_XI5/MM911_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1264 XI5/NET05362 N_NET29_XI5/MM1264_g N_VSS_XI5/MM1264_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM880 N_NET147_XI5/MM880_d N_NET30_XI5/MM880_g N_VSS_XI5/MM880_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1256 XI5/NET05318 N_NET31_XI5/MM1256_g N_VSS_XI5/MM1256_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM879 N_NET147_XI5/MM879_d N_NET32_XI5/MM879_g N_VSS_XI5/MM879_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1248 XI5/NET05286 N_NET33_XI5/MM1248_g N_VSS_XI5/MM1248_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM848 N_NET147_XI5/MM848_d N_NET34_XI5/MM848_g N_VSS_XI5/MM848_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1240 XI5/NET05254 N_NET35_XI5/MM1240_g N_VSS_XI5/MM1240_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM847 N_NET147_XI5/MM847_d N_NET36_XI5/MM847_g N_VSS_XI5/MM847_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1232 XI5/NET05222 N_NET37_XI5/MM1232_g N_VSS_XI5/MM1232_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM816 N_NET147_XI5/MM816_d N_NET38_XI5/MM816_g N_VSS_XI5/MM816_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1224 XI5/NET05182 N_NET39_XI5/MM1224_g N_VSS_XI5/MM1224_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM815 N_NET147_XI5/MM815_d N_NET40_XI5/MM815_g N_VSS_XI5/MM815_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1216 XI5/NET05150 N_NET41_XI5/MM1216_g N_VSS_XI5/MM1216_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM784 N_NET147_XI5/MM784_d N_NET42_XI5/MM784_g N_VSS_XI5/MM784_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1208 XI5/NET05114 N_NET43_XI5/MM1208_g N_VSS_XI5/MM1208_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM783 N_NET147_XI5/MM783_d N_NET44_XI5/MM783_g N_VSS_XI5/MM783_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1200 XI5/NET05082 N_NET45_XI5/MM1200_g N_VSS_XI5/MM1200_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM752 N_NET147_XI5/MM752_d N_NET46_XI5/MM752_g N_VSS_XI5/MM752_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1192 XI5/NET05050 N_NET47_XI5/MM1192_g N_VSS_XI5/MM1192_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM751 N_NET147_XI5/MM751_d N_NET48_XI5/MM751_g N_VSS_XI5/MM751_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1184 XI5/NET05018 N_NET49_XI5/MM1184_g N_VSS_XI5/MM1184_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM735 N_NET147_XI5/MM735_d N_NET50_XI5/MM735_g N_VSS_XI5/MM735_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1176 XI5/NET04986 N_NET51_XI5/MM1176_g N_VSS_XI5/MM1176_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM704 N_NET147_XI5/MM704_d N_NET52_XI5/MM704_g N_VSS_XI5/MM704_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1168 XI5/NET04954 N_NET53_XI5/MM1168_g N_VSS_XI5/MM1168_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM703 N_NET147_XI5/MM703_d N_NET54_XI5/MM703_g N_VSS_XI5/MM703_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1160 XI5/NET04914 N_NET55_XI5/MM1160_g N_VSS_XI5/MM1160_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM672 N_NET147_XI5/MM672_d N_NET56_XI5/MM672_g N_VSS_XI5/MM672_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1152 XI5/NET04882 N_NET57_XI5/MM1152_g N_VSS_XI5/MM1152_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM671 N_NET147_XI5/MM671_d N_NET58_XI5/MM671_g N_VSS_XI5/MM671_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1144 XI5/NET04850 N_NET59_XI5/MM1144_g N_VSS_XI5/MM1144_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM640 N_NET147_XI5/MM640_d N_NET60_XI5/MM640_g N_VSS_XI5/MM640_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1136 XI5/NET04818 N_NET61_XI5/MM1136_g N_VSS_XI5/MM1136_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM639 N_NET147_XI5/MM639_d N_NET62_XI5/MM639_g N_VSS_XI5/MM639_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1128 XI5/NET04766 N_NET63_XI5/MM1128_g N_VSS_XI5/MM1128_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM608 N_NET147_XI5/MM608_d N_NET64_XI5/MM608_g N_VSS_XI5/MM608_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1111 XI5/NET04734 N_NET65_XI5/MM1111_g N_VSS_XI5/MM1111_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM605 N_NET147_XI5/MM605_d N_NET66_XI5/MM605_g N_VSS_XI5/MM605_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1095 XI5/NET04654 N_NET67_XI5/MM1095_g N_VSS_XI5/MM1095_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM578 N_NET147_XI5/MM578_d N_NET68_XI5/MM578_g N_VSS_XI5/MM578_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1087 XI5/NET04618 N_NET69_XI5/MM1087_g N_VSS_XI5/MM1087_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM530 N_NET147_XI5/MM530_d N_NET70_XI5/MM530_g N_VSS_XI5/MM530_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1079 XI5/NET04586 N_NET71_XI5/MM1079_g N_VSS_XI5/MM1079_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM529 N_NET147_XI5/MM529_d N_NET72_XI5/MM529_g N_VSS_XI5/MM529_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1063 XI5/NET04390 N_NET8_XI5/MM1063_g N_VSS_XI5/MM1063_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM2 N_NET148_XI7/MM2_d N_XI7/NET48_XI7/MM2_g N_XI7/NET141_XI7/MM2_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI5/MM1585 XI5/NET01346 N_NET10_XI5/MM1585_g N_VSS_XI5/MM1585_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1041 N_NET148_XI5/MM1041_d N_NET11_XI5/MM1041_g N_VSS_XI5/MM1041_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1577 XI5/NET01378 N_NET12_XI5/MM1577_g N_VSS_XI5/MM1577_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1038 N_NET148_XI5/MM1038_d N_NET13_XI5/MM1038_g N_VSS_XI5/MM1038_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1569 XI5/NET01410 N_NET14_XI5/MM1569_g N_VSS_XI5/MM1569_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1009 N_NET148_XI5/MM1009_d N_NET15_XI5/MM1009_g N_VSS_XI5/MM1009_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1561 XI5/NET01442 N_NET16_XI5/MM1561_g N_VSS_XI5/MM1561_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1006 N_NET148_XI5/MM1006_d N_NET17_XI5/MM1006_g N_VSS_XI5/MM1006_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1553 XI5/NET01474 N_NET18_XI5/MM1553_g N_VSS_XI5/MM1553_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM977 N_NET148_XI5/MM977_d N_NET19_XI5/MM977_g N_VSS_XI5/MM977_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1545 XI5/NET01506 N_NET20_XI5/MM1545_g N_VSS_XI5/MM1545_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM974 N_NET148_XI5/MM974_d N_NET21_XI5/MM974_g N_VSS_XI5/MM974_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1537 XI5/NET01538 N_NET22_XI5/MM1537_g N_VSS_XI5/MM1537_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM945 N_NET148_XI5/MM945_d N_NET23_XI5/MM945_g N_VSS_XI5/MM945_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1529 XI5/NET01570 N_NET24_XI5/MM1529_g N_VSS_XI5/MM1529_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM942 N_NET148_XI5/MM942_d N_NET25_XI5/MM942_g N_VSS_XI5/MM942_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1521 XI5/NET01602 N_NET26_XI5/MM1521_g N_VSS_XI5/MM1521_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM913 N_NET148_XI5/MM913_d N_NET27_XI5/MM913_g N_VSS_XI5/MM913_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1513 XI5/NET01634 N_NET28_XI5/MM1513_g N_VSS_XI5/MM1513_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM910 N_NET148_XI5/MM910_d N_NET29_XI5/MM910_g N_VSS_XI5/MM910_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1505 XI5/NET01666 N_NET30_XI5/MM1505_g N_VSS_XI5/MM1505_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM881 N_NET148_XI5/MM881_d N_NET31_XI5/MM881_g N_VSS_XI5/MM881_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1497 XI5/NET01698 N_NET32_XI5/MM1497_g N_VSS_XI5/MM1497_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM878 N_NET148_XI5/MM878_d N_NET33_XI5/MM878_g N_VSS_XI5/MM878_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1489 XI5/NET01730 N_NET34_XI5/MM1489_g N_VSS_XI5/MM1489_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM849 N_NET148_XI5/MM849_d N_NET35_XI5/MM849_g N_VSS_XI5/MM849_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1481 XI5/NET01762 N_NET36_XI5/MM1481_g N_VSS_XI5/MM1481_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM846 N_NET148_XI5/MM846_d N_NET37_XI5/MM846_g N_VSS_XI5/MM846_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1473 XI5/NET01794 N_NET38_XI5/MM1473_g N_VSS_XI5/MM1473_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM817 N_NET148_XI5/MM817_d N_NET39_XI5/MM817_g N_VSS_XI5/MM817_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1465 XI5/NET01826 N_NET40_XI5/MM1465_g N_VSS_XI5/MM1465_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM814 N_NET148_XI5/MM814_d N_NET41_XI5/MM814_g N_VSS_XI5/MM814_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1457 XI5/NET01858 N_NET42_XI5/MM1457_g N_VSS_XI5/MM1457_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM785 N_NET148_XI5/MM785_d N_NET43_XI5/MM785_g N_VSS_XI5/MM785_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1449 XI5/NET01890 N_NET44_XI5/MM1449_g N_VSS_XI5/MM1449_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM782 N_NET148_XI5/MM782_d N_NET45_XI5/MM782_g N_VSS_XI5/MM782_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1441 XI5/NET01922 N_NET46_XI5/MM1441_g N_VSS_XI5/MM1441_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM753 N_NET148_XI5/MM753_d N_NET47_XI5/MM753_g N_VSS_XI5/MM753_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1433 XI5/NET01954 N_NET48_XI5/MM1433_g N_VSS_XI5/MM1433_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM750 N_NET148_XI5/MM750_d N_NET49_XI5/MM750_g N_VSS_XI5/MM750_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1425 XI5/NET01986 N_NET50_XI5/MM1425_g N_VSS_XI5/MM1425_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM734 N_NET148_XI5/MM734_d N_NET51_XI5/MM734_g N_VSS_XI5/MM734_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1417 XI5/NET02018 N_NET52_XI5/MM1417_g N_VSS_XI5/MM1417_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM705 N_NET148_XI5/MM705_d N_NET53_XI5/MM705_g N_VSS_XI5/MM705_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1409 XI5/NET02050 N_NET54_XI5/MM1409_g N_VSS_XI5/MM1409_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM702 N_NET148_XI5/MM702_d N_NET55_XI5/MM702_g N_VSS_XI5/MM702_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1401 XI5/NET02082 N_NET56_XI5/MM1401_g N_VSS_XI5/MM1401_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM673 N_NET148_XI5/MM673_d N_NET57_XI5/MM673_g N_VSS_XI5/MM673_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1393 XI5/NET02114 N_NET58_XI5/MM1393_g N_VSS_XI5/MM1393_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM670 N_NET148_XI5/MM670_d N_NET59_XI5/MM670_g N_VSS_XI5/MM670_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1385 XI5/NET02146 N_NET60_XI5/MM1385_g N_VSS_XI5/MM1385_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM641 N_NET148_XI5/MM641_d N_NET61_XI5/MM641_g N_VSS_XI5/MM641_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1377 XI5/NET02178 N_NET62_XI5/MM1377_g N_VSS_XI5/MM1377_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM638 N_NET148_XI5/MM638_d N_NET63_XI5/MM638_g N_VSS_XI5/MM638_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1369 XI5/NET02210 N_NET64_XI5/MM1369_g N_VSS_XI5/MM1369_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM609 N_NET148_XI5/MM609_d N_NET65_XI5/MM609_g N_VSS_XI5/MM609_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1361 XI5/NET02242 N_NET66_XI5/MM1361_g N_VSS_XI5/MM1361_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM592 N_NET148_XI5/MM592_d N_NET67_XI5/MM592_g N_VSS_XI5/MM592_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1353 XI5/NET02274 N_NET68_XI5/MM1353_g N_VSS_XI5/MM1353_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM591 N_NET148_XI5/MM591_d N_NET69_XI5/MM591_g N_VSS_XI5/MM591_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1352 XI5/NET02278 N_NET70_XI5/MM1352_g N_VSS_XI5/MM1352_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM545 N_NET148_XI5/MM545_d N_NET71_XI5/MM545_g N_VSS_XI5/MM545_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1071 XI5/NET04538 N_NET72_XI5/MM1071_g N_VSS_XI5/MM1071_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM0 N_NET148_XI5/MM0_d N_NET8_XI5/MM0_g N_VSS_XI5/MM0_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM23 N_XI7/NET141_XI7/MM23_d N_NET125_XI7/MM23_g N_XI7/NET101_XI7/MM23_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI7/MM22 N_XI7/NET125_XI7/MM22_d N_XI7/NET68_XI7/MM22_g N_XI7/NET101_XI7/MM22_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI7/MM11 N_NET149_XI7/MM11_d N_NET120_XI7/MM11_g N_XI7/NET125_XI7/MM11_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI5/MM1055 N_NET149_XI5/MM1055_d N_NET10_XI5/MM1055_g N_VSS_XI5/MM1055_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1336 XI5/NET02310 N_NET11_XI5/MM1336_g N_VSS_XI5/MM1336_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1024 N_NET149_XI5/MM1024_d N_NET12_XI5/MM1024_g N_VSS_XI5/MM1024_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1322 XI5/NET02366 N_NET13_XI5/MM1322_g N_VSS_XI5/MM1322_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1023 N_NET149_XI5/MM1023_d N_NET14_XI5/MM1023_g N_VSS_XI5/MM1023_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1314 XI5/NET02398 N_NET15_XI5/MM1314_g N_VSS_XI5/MM1314_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM992 N_NET149_XI5/MM992_d N_NET16_XI5/MM992_g N_VSS_XI5/MM992_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1306 XI5/NET02430 N_NET17_XI5/MM1306_g N_VSS_XI5/MM1306_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM991 N_NET149_XI5/MM991_d N_NET18_XI5/MM991_g N_VSS_XI5/MM991_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1298 XI5/NET02462 N_NET19_XI5/MM1298_g N_VSS_XI5/MM1298_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM960 N_NET149_XI5/MM960_d N_NET20_XI5/MM960_g N_VSS_XI5/MM960_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1290 XI5/NET04282 N_NET21_XI5/MM1290_g N_VSS_XI5/MM1290_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM959 N_NET149_XI5/MM959_d N_NET22_XI5/MM959_g N_VSS_XI5/MM959_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1282 XI5/NET04314 N_NET23_XI5/MM1282_g N_VSS_XI5/MM1282_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM928 N_NET149_XI5/MM928_d N_NET24_XI5/MM928_g N_VSS_XI5/MM928_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1274 XI5/NET03462 N_NET25_XI5/MM1274_g N_VSS_XI5/MM1274_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM927 N_NET149_XI5/MM927_d N_NET26_XI5/MM927_g N_VSS_XI5/MM927_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1271 XI5/NET05402 N_NET27_XI5/MM1271_g N_VSS_XI5/MM1271_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM896 N_NET149_XI5/MM896_d N_NET28_XI5/MM896_g N_VSS_XI5/MM896_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1263 XI5/NET05358 N_NET29_XI5/MM1263_g N_VSS_XI5/MM1263_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM895 N_NET149_XI5/MM895_d N_NET30_XI5/MM895_g N_VSS_XI5/MM895_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1255 XI5/NET05314 N_NET31_XI5/MM1255_g N_VSS_XI5/MM1255_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM864 N_NET149_XI5/MM864_d N_NET32_XI5/MM864_g N_VSS_XI5/MM864_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1247 XI5/NET05282 N_NET33_XI5/MM1247_g N_VSS_XI5/MM1247_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM863 N_NET149_XI5/MM863_d N_NET34_XI5/MM863_g N_VSS_XI5/MM863_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1239 XI5/NET05250 N_NET35_XI5/MM1239_g N_VSS_XI5/MM1239_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM832 N_NET149_XI5/MM832_d N_NET36_XI5/MM832_g N_VSS_XI5/MM832_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1231 XI5/NET05218 N_NET37_XI5/MM1231_g N_VSS_XI5/MM1231_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM831 N_NET149_XI5/MM831_d N_NET38_XI5/MM831_g N_VSS_XI5/MM831_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1223 XI5/NET05178 N_NET39_XI5/MM1223_g N_VSS_XI5/MM1223_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM800 N_NET149_XI5/MM800_d N_NET40_XI5/MM800_g N_VSS_XI5/MM800_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1215 XI5/NET05146 N_NET41_XI5/MM1215_g N_VSS_XI5/MM1215_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM799 N_NET149_XI5/MM799_d N_NET42_XI5/MM799_g N_VSS_XI5/MM799_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1207 XI5/NET05110 N_NET43_XI5/MM1207_g N_VSS_XI5/MM1207_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM768 N_NET149_XI5/MM768_d N_NET44_XI5/MM768_g N_VSS_XI5/MM768_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1199 XI5/NET05078 N_NET45_XI5/MM1199_g N_VSS_XI5/MM1199_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM767 N_NET149_XI5/MM767_d N_NET46_XI5/MM767_g N_VSS_XI5/MM767_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1191 XI5/NET05046 N_NET47_XI5/MM1191_g N_VSS_XI5/MM1191_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM736 N_NET149_XI5/MM736_d N_NET48_XI5/MM736_g N_VSS_XI5/MM736_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1183 XI5/NET05014 N_NET49_XI5/MM1183_g N_VSS_XI5/MM1183_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM720 N_NET149_XI5/MM720_d N_NET50_XI5/MM720_g N_VSS_XI5/MM720_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1175 XI5/NET04982 N_NET51_XI5/MM1175_g N_VSS_XI5/MM1175_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM719 N_NET149_XI5/MM719_d N_NET52_XI5/MM719_g N_VSS_XI5/MM719_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1167 XI5/NET04950 N_NET53_XI5/MM1167_g N_VSS_XI5/MM1167_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM688 N_NET149_XI5/MM688_d N_NET54_XI5/MM688_g N_VSS_XI5/MM688_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1159 XI5/NET04910 N_NET55_XI5/MM1159_g N_VSS_XI5/MM1159_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM687 N_NET149_XI5/MM687_d N_NET56_XI5/MM687_g N_VSS_XI5/MM687_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1151 XI5/NET04878 N_NET57_XI5/MM1151_g N_VSS_XI5/MM1151_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM656 N_NET149_XI5/MM656_d N_NET58_XI5/MM656_g N_VSS_XI5/MM656_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1143 XI5/NET04846 N_NET59_XI5/MM1143_g N_VSS_XI5/MM1143_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM655 N_NET149_XI5/MM655_d N_NET60_XI5/MM655_g N_VSS_XI5/MM655_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1135 XI5/NET04814 N_NET61_XI5/MM1135_g N_VSS_XI5/MM1135_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM624 N_NET149_XI5/MM624_d N_NET62_XI5/MM624_g N_VSS_XI5/MM624_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1127 XI5/NET04762 N_NET63_XI5/MM1127_g N_VSS_XI5/MM1127_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM623 N_NET149_XI5/MM623_d N_NET64_XI5/MM623_g N_VSS_XI5/MM623_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1110 XI5/NET04730 N_NET65_XI5/MM1110_g N_VSS_XI5/MM1110_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM607 N_NET149_XI5/MM607_d N_NET66_XI5/MM607_g N_VSS_XI5/MM607_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1094 XI5/NET04650 N_NET67_XI5/MM1094_g N_VSS_XI5/MM1094_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM576 N_NET149_XI5/MM576_d N_NET68_XI5/MM576_g N_VSS_XI5/MM576_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1086 XI5/NET04614 N_NET69_XI5/MM1086_g N_VSS_XI5/MM1086_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM535 N_NET149_XI5/MM535_d N_NET70_XI5/MM535_g N_VSS_XI5/MM535_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1078 XI5/NET04582 N_NET71_XI5/MM1078_g N_VSS_XI5/MM1078_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM524 N_NET149_XI5/MM524_d N_NET72_XI5/MM524_g N_VSS_XI5/MM524_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1062 XI5/NET04386 N_NET8_XI5/MM1062_g N_VSS_XI5/MM1062_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM10 N_NET151_XI7/MM10_d N_XI7/NET48_XI7/MM10_g N_XI7/NET125_XI7/MM10_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI5/MM1586 XI5/NET01342 N_NET10_XI5/MM1586_g N_VSS_XI5/MM1586_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1046 N_NET151_XI5/MM1046_d N_NET11_XI5/MM1046_g N_VSS_XI5/MM1046_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1578 XI5/NET01374 N_NET12_XI5/MM1578_g N_VSS_XI5/MM1578_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1033 N_NET151_XI5/MM1033_d N_NET13_XI5/MM1033_g N_VSS_XI5/MM1033_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1570 XI5/NET01406 N_NET14_XI5/MM1570_g N_VSS_XI5/MM1570_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1014 N_NET151_XI5/MM1014_d N_NET15_XI5/MM1014_g N_VSS_XI5/MM1014_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1562 XI5/NET01438 N_NET16_XI5/MM1562_g N_VSS_XI5/MM1562_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1001 N_NET151_XI5/MM1001_d N_NET17_XI5/MM1001_g N_VSS_XI5/MM1001_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1554 XI5/NET01470 N_NET18_XI5/MM1554_g N_VSS_XI5/MM1554_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM982 N_NET151_XI5/MM982_d N_NET19_XI5/MM982_g N_VSS_XI5/MM982_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1546 XI5/NET01502 N_NET20_XI5/MM1546_g N_VSS_XI5/MM1546_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM969 N_NET151_XI5/MM969_d N_NET21_XI5/MM969_g N_VSS_XI5/MM969_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1538 XI5/NET01534 N_NET22_XI5/MM1538_g N_VSS_XI5/MM1538_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM950 N_NET151_XI5/MM950_d N_NET23_XI5/MM950_g N_VSS_XI5/MM950_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1530 XI5/NET01566 N_NET24_XI5/MM1530_g N_VSS_XI5/MM1530_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM937 N_NET151_XI5/MM937_d N_NET25_XI5/MM937_g N_VSS_XI5/MM937_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1522 XI5/NET01598 N_NET26_XI5/MM1522_g N_VSS_XI5/MM1522_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM918 N_NET151_XI5/MM918_d N_NET27_XI5/MM918_g N_VSS_XI5/MM918_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1514 XI5/NET01630 N_NET28_XI5/MM1514_g N_VSS_XI5/MM1514_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM905 N_NET151_XI5/MM905_d N_NET29_XI5/MM905_g N_VSS_XI5/MM905_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1506 XI5/NET01662 N_NET30_XI5/MM1506_g N_VSS_XI5/MM1506_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM886 N_NET151_XI5/MM886_d N_NET31_XI5/MM886_g N_VSS_XI5/MM886_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1498 XI5/NET01694 N_NET32_XI5/MM1498_g N_VSS_XI5/MM1498_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM873 N_NET151_XI5/MM873_d N_NET33_XI5/MM873_g N_VSS_XI5/MM873_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1490 XI5/NET01726 N_NET34_XI5/MM1490_g N_VSS_XI5/MM1490_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM854 N_NET151_XI5/MM854_d N_NET35_XI5/MM854_g N_VSS_XI5/MM854_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1482 XI5/NET01758 N_NET36_XI5/MM1482_g N_VSS_XI5/MM1482_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM841 N_NET151_XI5/MM841_d N_NET37_XI5/MM841_g N_VSS_XI5/MM841_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1474 XI5/NET01790 N_NET38_XI5/MM1474_g N_VSS_XI5/MM1474_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM822 N_NET151_XI5/MM822_d N_NET39_XI5/MM822_g N_VSS_XI5/MM822_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1466 XI5/NET01822 N_NET40_XI5/MM1466_g N_VSS_XI5/MM1466_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM809 N_NET151_XI5/MM809_d N_NET41_XI5/MM809_g N_VSS_XI5/MM809_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1458 XI5/NET01854 N_NET42_XI5/MM1458_g N_VSS_XI5/MM1458_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM790 N_NET151_XI5/MM790_d N_NET43_XI5/MM790_g N_VSS_XI5/MM790_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1450 XI5/NET01886 N_NET44_XI5/MM1450_g N_VSS_XI5/MM1450_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM777 N_NET151_XI5/MM777_d N_NET45_XI5/MM777_g N_VSS_XI5/MM777_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1442 XI5/NET01918 N_NET46_XI5/MM1442_g N_VSS_XI5/MM1442_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM758 N_NET151_XI5/MM758_d N_NET47_XI5/MM758_g N_VSS_XI5/MM758_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1434 XI5/NET01950 N_NET48_XI5/MM1434_g N_VSS_XI5/MM1434_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM745 N_NET151_XI5/MM745_d N_NET49_XI5/MM745_g N_VSS_XI5/MM745_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1426 XI5/NET01982 N_NET50_XI5/MM1426_g N_VSS_XI5/MM1426_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM729 N_NET151_XI5/MM729_d N_NET51_XI5/MM729_g N_VSS_XI5/MM729_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1418 XI5/NET02014 N_NET52_XI5/MM1418_g N_VSS_XI5/MM1418_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM710 N_NET151_XI5/MM710_d N_NET53_XI5/MM710_g N_VSS_XI5/MM710_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1410 XI5/NET02046 N_NET54_XI5/MM1410_g N_VSS_XI5/MM1410_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM697 N_NET151_XI5/MM697_d N_NET55_XI5/MM697_g N_VSS_XI5/MM697_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1402 XI5/NET02078 N_NET56_XI5/MM1402_g N_VSS_XI5/MM1402_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM678 N_NET151_XI5/MM678_d N_NET57_XI5/MM678_g N_VSS_XI5/MM678_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1394 XI5/NET02110 N_NET58_XI5/MM1394_g N_VSS_XI5/MM1394_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM665 N_NET151_XI5/MM665_d N_NET59_XI5/MM665_g N_VSS_XI5/MM665_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1386 XI5/NET02142 N_NET60_XI5/MM1386_g N_VSS_XI5/MM1386_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM646 N_NET151_XI5/MM646_d N_NET61_XI5/MM646_g N_VSS_XI5/MM646_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1378 XI5/NET02174 N_NET62_XI5/MM1378_g N_VSS_XI5/MM1378_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM633 N_NET151_XI5/MM633_d N_NET63_XI5/MM633_g N_VSS_XI5/MM633_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1370 XI5/NET02206 N_NET64_XI5/MM1370_g N_VSS_XI5/MM1370_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM614 N_NET151_XI5/MM614_d N_NET65_XI5/MM614_g N_VSS_XI5/MM614_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1362 XI5/NET02238 N_NET66_XI5/MM1362_g N_VSS_XI5/MM1362_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM597 N_NET151_XI5/MM597_d N_NET67_XI5/MM597_g N_VSS_XI5/MM597_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1354 XI5/NET02270 N_NET68_XI5/MM1354_g N_VSS_XI5/MM1354_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM586 N_NET151_XI5/MM586_d N_NET69_XI5/MM586_g N_VSS_XI5/MM586_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1351 XI5/NET02282 N_NET70_XI5/MM1351_g N_VSS_XI5/MM1351_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM540 N_NET151_XI5/MM540_d N_NET71_XI5/MM540_g N_VSS_XI5/MM540_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1070 XI5/NET04534 N_NET72_XI5/MM1070_g N_VSS_XI5/MM1070_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM515 N_NET151_XI5/MM515_d N_NET8_XI5/MM515_g N_VSS_XI5/MM515_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM30 N_XI7/NET101_XI7/MM30_d N_NET85_XI7/MM30_g N_NET139_XI7/MM30_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI7/MM31 N_XI7/NET89_XI7/MM31_d N_XI7/NET76_XI7/MM31_g N_NET139_XI7/MM31_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI7/MM16 N_NET152_XI7/MM16_d N_NET120_XI7/MM16_g N_XI7/NET113_XI7/MM16_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI5/MM1053 N_NET152_XI5/MM1053_d N_NET10_XI5/MM1053_g N_VSS_XI5/MM1053_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1329 XI5/NET02338 N_NET11_XI5/MM1329_g N_VSS_XI5/MM1329_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1026 N_NET152_XI5/MM1026_d N_NET12_XI5/MM1026_g N_VSS_XI5/MM1026_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1323 XI5/NET02362 N_NET13_XI5/MM1323_g N_VSS_XI5/MM1323_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1021 N_NET152_XI5/MM1021_d N_NET14_XI5/MM1021_g N_VSS_XI5/MM1021_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1315 XI5/NET02394 N_NET15_XI5/MM1315_g N_VSS_XI5/MM1315_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM994 N_NET152_XI5/MM994_d N_NET16_XI5/MM994_g N_VSS_XI5/MM994_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1307 XI5/NET02426 N_NET17_XI5/MM1307_g N_VSS_XI5/MM1307_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM989 N_NET152_XI5/MM989_d N_NET18_XI5/MM989_g N_VSS_XI5/MM989_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1299 XI5/NET02458 N_NET19_XI5/MM1299_g N_VSS_XI5/MM1299_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM962 N_NET152_XI5/MM962_d N_NET20_XI5/MM962_g N_VSS_XI5/MM962_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1291 XI5/NET04278 N_NET21_XI5/MM1291_g N_VSS_XI5/MM1291_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM957 N_NET152_XI5/MM957_d N_NET22_XI5/MM957_g N_VSS_XI5/MM957_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1283 XI5/NET04310 N_NET23_XI5/MM1283_g N_VSS_XI5/MM1283_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM930 N_NET152_XI5/MM930_d N_NET24_XI5/MM930_g N_VSS_XI5/MM930_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1275 XI5/NET03458 N_NET25_XI5/MM1275_g N_VSS_XI5/MM1275_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM925 N_NET152_XI5/MM925_d N_NET26_XI5/MM925_g N_VSS_XI5/MM925_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1270 XI5/NET05398 N_NET27_XI5/MM1270_g N_VSS_XI5/MM1270_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM898 N_NET152_XI5/MM898_d N_NET28_XI5/MM898_g N_VSS_XI5/MM898_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1262 XI5/NET05354 N_NET29_XI5/MM1262_g N_VSS_XI5/MM1262_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM893 N_NET152_XI5/MM893_d N_NET30_XI5/MM893_g N_VSS_XI5/MM893_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1254 XI5/NET05310 N_NET31_XI5/MM1254_g N_VSS_XI5/MM1254_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM866 N_NET152_XI5/MM866_d N_NET32_XI5/MM866_g N_VSS_XI5/MM866_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1246 XI5/NET05278 N_NET33_XI5/MM1246_g N_VSS_XI5/MM1246_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM861 N_NET152_XI5/MM861_d N_NET34_XI5/MM861_g N_VSS_XI5/MM861_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1238 XI5/NET05246 N_NET35_XI5/MM1238_g N_VSS_XI5/MM1238_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM834 N_NET152_XI5/MM834_d N_NET36_XI5/MM834_g N_VSS_XI5/MM834_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1230 XI5/NET05214 N_NET37_XI5/MM1230_g N_VSS_XI5/MM1230_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM829 N_NET152_XI5/MM829_d N_NET38_XI5/MM829_g N_VSS_XI5/MM829_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1222 XI5/NET05174 N_NET39_XI5/MM1222_g N_VSS_XI5/MM1222_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM802 N_NET152_XI5/MM802_d N_NET40_XI5/MM802_g N_VSS_XI5/MM802_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1214 XI5/NET05142 N_NET41_XI5/MM1214_g N_VSS_XI5/MM1214_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM797 N_NET152_XI5/MM797_d N_NET42_XI5/MM797_g N_VSS_XI5/MM797_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1206 XI5/NET05106 N_NET43_XI5/MM1206_g N_VSS_XI5/MM1206_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM770 N_NET152_XI5/MM770_d N_NET44_XI5/MM770_g N_VSS_XI5/MM770_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1198 XI5/NET05074 N_NET45_XI5/MM1198_g N_VSS_XI5/MM1198_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM765 N_NET152_XI5/MM765_d N_NET46_XI5/MM765_g N_VSS_XI5/MM765_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1190 XI5/NET05042 N_NET47_XI5/MM1190_g N_VSS_XI5/MM1190_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM738 N_NET152_XI5/MM738_d N_NET48_XI5/MM738_g N_VSS_XI5/MM738_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1182 XI5/NET05010 N_NET49_XI5/MM1182_g N_VSS_XI5/MM1182_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM722 N_NET152_XI5/MM722_d N_NET50_XI5/MM722_g N_VSS_XI5/MM722_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1174 XI5/NET04978 N_NET51_XI5/MM1174_g N_VSS_XI5/MM1174_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM717 N_NET152_XI5/MM717_d N_NET52_XI5/MM717_g N_VSS_XI5/MM717_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1166 XI5/NET04946 N_NET53_XI5/MM1166_g N_VSS_XI5/MM1166_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM690 N_NET152_XI5/MM690_d N_NET54_XI5/MM690_g N_VSS_XI5/MM690_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1158 XI5/NET04906 N_NET55_XI5/MM1158_g N_VSS_XI5/MM1158_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM685 N_NET152_XI5/MM685_d N_NET56_XI5/MM685_g N_VSS_XI5/MM685_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1150 XI5/NET04874 N_NET57_XI5/MM1150_g N_VSS_XI5/MM1150_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM658 N_NET152_XI5/MM658_d N_NET58_XI5/MM658_g N_VSS_XI5/MM658_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1142 XI5/NET04842 N_NET59_XI5/MM1142_g N_VSS_XI5/MM1142_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM653 N_NET152_XI5/MM653_d N_NET60_XI5/MM653_g N_VSS_XI5/MM653_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1134 XI5/NET04810 N_NET61_XI5/MM1134_g N_VSS_XI5/MM1134_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM626 N_NET152_XI5/MM626_d N_NET62_XI5/MM626_g N_VSS_XI5/MM626_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1126 XI5/NET04758 N_NET63_XI5/MM1126_g N_VSS_XI5/MM1126_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM621 N_NET152_XI5/MM621_d N_NET64_XI5/MM621_g N_VSS_XI5/MM621_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1109 XI5/NET04722 N_NET65_XI5/MM1109_g N_VSS_XI5/MM1109_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM604 N_NET152_XI5/MM604_d N_NET66_XI5/MM604_g N_VSS_XI5/MM604_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1093 XI5/NET04642 N_NET67_XI5/MM1093_g N_VSS_XI5/MM1093_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM579 N_NET152_XI5/MM579_d N_NET68_XI5/MM579_g N_VSS_XI5/MM579_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1085 XI5/NET04610 N_NET69_XI5/MM1085_g N_VSS_XI5/MM1085_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM533 N_NET152_XI5/MM533_d N_NET70_XI5/MM533_g N_VSS_XI5/MM533_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1077 XI5/NET04578 N_NET71_XI5/MM1077_g N_VSS_XI5/MM1077_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM526 N_NET152_XI5/MM526_d N_NET72_XI5/MM526_g N_VSS_XI5/MM526_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1061 XI5/NET04382 N_NET8_XI5/MM1061_g N_VSS_XI5/MM1061_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM17 N_NET153_XI7/MM17_d N_XI7/NET48_XI7/MM17_g N_XI7/NET113_XI7/MM17_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI5/MM1587 XI5/NET01338 N_NET10_XI5/MM1587_g N_VSS_XI5/MM1587_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1044 N_NET153_XI5/MM1044_d N_NET11_XI5/MM1044_g N_VSS_XI5/MM1044_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1579 XI5/NET01370 N_NET12_XI5/MM1579_g N_VSS_XI5/MM1579_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1035 N_NET153_XI5/MM1035_d N_NET13_XI5/MM1035_g N_VSS_XI5/MM1035_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1571 XI5/NET01402 N_NET14_XI5/MM1571_g N_VSS_XI5/MM1571_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1012 N_NET153_XI5/MM1012_d N_NET15_XI5/MM1012_g N_VSS_XI5/MM1012_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1563 XI5/NET01434 N_NET16_XI5/MM1563_g N_VSS_XI5/MM1563_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1003 N_NET153_XI5/MM1003_d N_NET17_XI5/MM1003_g N_VSS_XI5/MM1003_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1555 XI5/NET01466 N_NET18_XI5/MM1555_g N_VSS_XI5/MM1555_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM980 N_NET153_XI5/MM980_d N_NET19_XI5/MM980_g N_VSS_XI5/MM980_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1547 XI5/NET01498 N_NET20_XI5/MM1547_g N_VSS_XI5/MM1547_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM971 N_NET153_XI5/MM971_d N_NET21_XI5/MM971_g N_VSS_XI5/MM971_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1539 XI5/NET01530 N_NET22_XI5/MM1539_g N_VSS_XI5/MM1539_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM948 N_NET153_XI5/MM948_d N_NET23_XI5/MM948_g N_VSS_XI5/MM948_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1531 XI5/NET01562 N_NET24_XI5/MM1531_g N_VSS_XI5/MM1531_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM939 N_NET153_XI5/MM939_d N_NET25_XI5/MM939_g N_VSS_XI5/MM939_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1523 XI5/NET01594 N_NET26_XI5/MM1523_g N_VSS_XI5/MM1523_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM916 N_NET153_XI5/MM916_d N_NET27_XI5/MM916_g N_VSS_XI5/MM916_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1515 XI5/NET01626 N_NET28_XI5/MM1515_g N_VSS_XI5/MM1515_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM907 N_NET153_XI5/MM907_d N_NET29_XI5/MM907_g N_VSS_XI5/MM907_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1507 XI5/NET01658 N_NET30_XI5/MM1507_g N_VSS_XI5/MM1507_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM884 N_NET153_XI5/MM884_d N_NET31_XI5/MM884_g N_VSS_XI5/MM884_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1499 XI5/NET01690 N_NET32_XI5/MM1499_g N_VSS_XI5/MM1499_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM875 N_NET153_XI5/MM875_d N_NET33_XI5/MM875_g N_VSS_XI5/MM875_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1491 XI5/NET01722 N_NET34_XI5/MM1491_g N_VSS_XI5/MM1491_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM852 N_NET153_XI5/MM852_d N_NET35_XI5/MM852_g N_VSS_XI5/MM852_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1483 XI5/NET01754 N_NET36_XI5/MM1483_g N_VSS_XI5/MM1483_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM843 N_NET153_XI5/MM843_d N_NET37_XI5/MM843_g N_VSS_XI5/MM843_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1475 XI5/NET01786 N_NET38_XI5/MM1475_g N_VSS_XI5/MM1475_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM820 N_NET153_XI5/MM820_d N_NET39_XI5/MM820_g N_VSS_XI5/MM820_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1467 XI5/NET01818 N_NET40_XI5/MM1467_g N_VSS_XI5/MM1467_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM811 N_NET153_XI5/MM811_d N_NET41_XI5/MM811_g N_VSS_XI5/MM811_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1459 XI5/NET01850 N_NET42_XI5/MM1459_g N_VSS_XI5/MM1459_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM788 N_NET153_XI5/MM788_d N_NET43_XI5/MM788_g N_VSS_XI5/MM788_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1451 XI5/NET01882 N_NET44_XI5/MM1451_g N_VSS_XI5/MM1451_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM779 N_NET153_XI5/MM779_d N_NET45_XI5/MM779_g N_VSS_XI5/MM779_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1443 XI5/NET01914 N_NET46_XI5/MM1443_g N_VSS_XI5/MM1443_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM756 N_NET153_XI5/MM756_d N_NET47_XI5/MM756_g N_VSS_XI5/MM756_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1435 XI5/NET01946 N_NET48_XI5/MM1435_g N_VSS_XI5/MM1435_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM747 N_NET153_XI5/MM747_d N_NET49_XI5/MM747_g N_VSS_XI5/MM747_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1427 XI5/NET01978 N_NET50_XI5/MM1427_g N_VSS_XI5/MM1427_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM731 N_NET153_XI5/MM731_d N_NET51_XI5/MM731_g N_VSS_XI5/MM731_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1419 XI5/NET02010 N_NET52_XI5/MM1419_g N_VSS_XI5/MM1419_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM708 N_NET153_XI5/MM708_d N_NET53_XI5/MM708_g N_VSS_XI5/MM708_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1411 XI5/NET02042 N_NET54_XI5/MM1411_g N_VSS_XI5/MM1411_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM699 N_NET153_XI5/MM699_d N_NET55_XI5/MM699_g N_VSS_XI5/MM699_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1403 XI5/NET02074 N_NET56_XI5/MM1403_g N_VSS_XI5/MM1403_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM676 N_NET153_XI5/MM676_d N_NET57_XI5/MM676_g N_VSS_XI5/MM676_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1395 XI5/NET02106 N_NET58_XI5/MM1395_g N_VSS_XI5/MM1395_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM667 N_NET153_XI5/MM667_d N_NET59_XI5/MM667_g N_VSS_XI5/MM667_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1387 XI5/NET02138 N_NET60_XI5/MM1387_g N_VSS_XI5/MM1387_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM644 N_NET153_XI5/MM644_d N_NET61_XI5/MM644_g N_VSS_XI5/MM644_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1379 XI5/NET02170 N_NET62_XI5/MM1379_g N_VSS_XI5/MM1379_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM635 N_NET153_XI5/MM635_d N_NET63_XI5/MM635_g N_VSS_XI5/MM635_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1371 XI5/NET02202 N_NET64_XI5/MM1371_g N_VSS_XI5/MM1371_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM612 N_NET153_XI5/MM612_d N_NET65_XI5/MM612_g N_VSS_XI5/MM612_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1363 XI5/NET02234 N_NET66_XI5/MM1363_g N_VSS_XI5/MM1363_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM595 N_NET153_XI5/MM595_d N_NET67_XI5/MM595_g N_VSS_XI5/MM595_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1355 XI5/NET02266 N_NET68_XI5/MM1355_g N_VSS_XI5/MM1355_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM588 N_NET153_XI5/MM588_d N_NET69_XI5/MM588_g N_VSS_XI5/MM588_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1349 XI5/NET02290 N_NET70_XI5/MM1349_g N_VSS_XI5/MM1349_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM542 N_NET153_XI5/MM542_d N_NET71_XI5/MM542_g N_VSS_XI5/MM542_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1069 XI5/NET04522 N_NET72_XI5/MM1069_g N_VSS_XI5/MM1069_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM517 N_NET153_XI5/MM517_d N_NET8_XI5/MM517_g N_VSS_XI5/MM517_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM26 N_XI7/NET113_XI7/MM26_d N_NET125_XI7/MM26_g N_XI7/NET89_XI7/MM26_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI7/MM27 N_XI7/NET109_XI7/MM27_d N_XI7/NET68_XI7/MM27_g N_XI7/NET89_XI7/MM27_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI7/MM19 N_NET154_XI7/MM19_d N_NET120_XI7/MM19_g N_XI7/NET109_XI7/MM19_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI5/MM1051 N_NET154_XI5/MM1051_d N_NET10_XI5/MM1051_g N_VSS_XI5/MM1051_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1333 XI5/NET02322 N_NET11_XI5/MM1333_g N_VSS_XI5/MM1333_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1028 N_NET154_XI5/MM1028_d N_NET12_XI5/MM1028_g N_VSS_XI5/MM1028_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1324 XI5/NET02358 N_NET13_XI5/MM1324_g N_VSS_XI5/MM1324_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1019 N_NET154_XI5/MM1019_d N_NET14_XI5/MM1019_g N_VSS_XI5/MM1019_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1316 XI5/NET02390 N_NET15_XI5/MM1316_g N_VSS_XI5/MM1316_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM996 N_NET154_XI5/MM996_d N_NET16_XI5/MM996_g N_VSS_XI5/MM996_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1308 XI5/NET02422 N_NET17_XI5/MM1308_g N_VSS_XI5/MM1308_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM987 N_NET154_XI5/MM987_d N_NET18_XI5/MM987_g N_VSS_XI5/MM987_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1300 XI5/NET02454 N_NET19_XI5/MM1300_g N_VSS_XI5/MM1300_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM964 N_NET154_XI5/MM964_d N_NET20_XI5/MM964_g N_VSS_XI5/MM964_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1292 XI5/NET04274 N_NET21_XI5/MM1292_g N_VSS_XI5/MM1292_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM955 N_NET154_XI5/MM955_d N_NET22_XI5/MM955_g N_VSS_XI5/MM955_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1284 XI5/NET04306 N_NET23_XI5/MM1284_g N_VSS_XI5/MM1284_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM932 N_NET154_XI5/MM932_d N_NET24_XI5/MM932_g N_VSS_XI5/MM932_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1276 XI5/NET03454 N_NET25_XI5/MM1276_g N_VSS_XI5/MM1276_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM923 N_NET154_XI5/MM923_d N_NET26_XI5/MM923_g N_VSS_XI5/MM923_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1269 XI5/NET05394 N_NET27_XI5/MM1269_g N_VSS_XI5/MM1269_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM900 N_NET154_XI5/MM900_d N_NET28_XI5/MM900_g N_VSS_XI5/MM900_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1261 XI5/NET05350 N_NET29_XI5/MM1261_g N_VSS_XI5/MM1261_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM891 N_NET154_XI5/MM891_d N_NET30_XI5/MM891_g N_VSS_XI5/MM891_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1253 XI5/NET05306 N_NET31_XI5/MM1253_g N_VSS_XI5/MM1253_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM868 N_NET154_XI5/MM868_d N_NET32_XI5/MM868_g N_VSS_XI5/MM868_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1245 XI5/NET05274 N_NET33_XI5/MM1245_g N_VSS_XI5/MM1245_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM859 N_NET154_XI5/MM859_d N_NET34_XI5/MM859_g N_VSS_XI5/MM859_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1237 XI5/NET05242 N_NET35_XI5/MM1237_g N_VSS_XI5/MM1237_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM836 N_NET154_XI5/MM836_d N_NET36_XI5/MM836_g N_VSS_XI5/MM836_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1229 XI5/NET05210 N_NET37_XI5/MM1229_g N_VSS_XI5/MM1229_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM827 N_NET154_XI5/MM827_d N_NET38_XI5/MM827_g N_VSS_XI5/MM827_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1221 XI5/NET05170 N_NET39_XI5/MM1221_g N_VSS_XI5/MM1221_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM804 N_NET154_XI5/MM804_d N_NET40_XI5/MM804_g N_VSS_XI5/MM804_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1213 XI5/NET05138 N_NET41_XI5/MM1213_g N_VSS_XI5/MM1213_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM795 N_NET154_XI5/MM795_d N_NET42_XI5/MM795_g N_VSS_XI5/MM795_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1205 XI5/NET05102 N_NET43_XI5/MM1205_g N_VSS_XI5/MM1205_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM772 N_NET154_XI5/MM772_d N_NET44_XI5/MM772_g N_VSS_XI5/MM772_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1197 XI5/NET05070 N_NET45_XI5/MM1197_g N_VSS_XI5/MM1197_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM763 N_NET154_XI5/MM763_d N_NET46_XI5/MM763_g N_VSS_XI5/MM763_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1189 XI5/NET05038 N_NET47_XI5/MM1189_g N_VSS_XI5/MM1189_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM740 N_NET154_XI5/MM740_d N_NET48_XI5/MM740_g N_VSS_XI5/MM740_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1181 XI5/NET05006 N_NET49_XI5/MM1181_g N_VSS_XI5/MM1181_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM724 N_NET154_XI5/MM724_d N_NET50_XI5/MM724_g N_VSS_XI5/MM724_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1173 XI5/NET04974 N_NET51_XI5/MM1173_g N_VSS_XI5/MM1173_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM715 N_NET154_XI5/MM715_d N_NET52_XI5/MM715_g N_VSS_XI5/MM715_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1165 XI5/NET04942 N_NET53_XI5/MM1165_g N_VSS_XI5/MM1165_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM692 N_NET154_XI5/MM692_d N_NET54_XI5/MM692_g N_VSS_XI5/MM692_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1157 XI5/NET04902 N_NET55_XI5/MM1157_g N_VSS_XI5/MM1157_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM683 N_NET154_XI5/MM683_d N_NET56_XI5/MM683_g N_VSS_XI5/MM683_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1149 XI5/NET04870 N_NET57_XI5/MM1149_g N_VSS_XI5/MM1149_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM660 N_NET154_XI5/MM660_d N_NET58_XI5/MM660_g N_VSS_XI5/MM660_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1141 XI5/NET04838 N_NET59_XI5/MM1141_g N_VSS_XI5/MM1141_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM651 N_NET154_XI5/MM651_d N_NET60_XI5/MM651_g N_VSS_XI5/MM651_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1133 XI5/NET04806 N_NET61_XI5/MM1133_g N_VSS_XI5/MM1133_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM628 N_NET154_XI5/MM628_d N_NET62_XI5/MM628_g N_VSS_XI5/MM628_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1125 XI5/NET04754 N_NET63_XI5/MM1125_g N_VSS_XI5/MM1125_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM619 N_NET154_XI5/MM619_d N_NET64_XI5/MM619_g N_VSS_XI5/MM619_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1108 XI5/NET04714 N_NET65_XI5/MM1108_g N_VSS_XI5/MM1108_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM602 N_NET154_XI5/MM602_d N_NET66_XI5/MM602_g N_VSS_XI5/MM602_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1092 XI5/NET04638 N_NET67_XI5/MM1092_g N_VSS_XI5/MM1092_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM581 N_NET154_XI5/MM581_d N_NET68_XI5/MM581_g N_VSS_XI5/MM581_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1084 XI5/NET04606 N_NET69_XI5/MM1084_g N_VSS_XI5/MM1084_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM536 N_NET154_XI5/MM536_d N_NET70_XI5/MM536_g N_VSS_XI5/MM536_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1076 XI5/NET04570 N_NET71_XI5/MM1076_g N_VSS_XI5/MM1076_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM523 N_NET154_XI5/MM523_d N_NET72_XI5/MM523_g N_VSS_XI5/MM523_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1060 XI5/NET04374 N_NET8_XI5/MM1060_g N_VSS_XI5/MM1060_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM18 N_NET155_XI7/MM18_d N_XI7/NET48_XI7/MM18_g N_XI7/NET109_XI7/MM18_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI5/MM1588 XI5/NET01334 N_NET10_XI5/MM1588_g N_VSS_XI5/MM1588_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1047 N_NET155_XI5/MM1047_d N_NET11_XI5/MM1047_g N_VSS_XI5/MM1047_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1580 XI5/NET01366 N_NET12_XI5/MM1580_g N_VSS_XI5/MM1580_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1032 N_NET155_XI5/MM1032_d N_NET13_XI5/MM1032_g N_VSS_XI5/MM1032_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1572 XI5/NET01398 N_NET14_XI5/MM1572_g N_VSS_XI5/MM1572_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1015 N_NET155_XI5/MM1015_d N_NET15_XI5/MM1015_g N_VSS_XI5/MM1015_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1564 XI5/NET01430 N_NET16_XI5/MM1564_g N_VSS_XI5/MM1564_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1000 N_NET155_XI5/MM1000_d N_NET17_XI5/MM1000_g N_VSS_XI5/MM1000_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1556 XI5/NET01462 N_NET18_XI5/MM1556_g N_VSS_XI5/MM1556_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM983 N_NET155_XI5/MM983_d N_NET19_XI5/MM983_g N_VSS_XI5/MM983_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1548 XI5/NET01494 N_NET20_XI5/MM1548_g N_VSS_XI5/MM1548_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM968 N_NET155_XI5/MM968_d N_NET21_XI5/MM968_g N_VSS_XI5/MM968_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1540 XI5/NET01526 N_NET22_XI5/MM1540_g N_VSS_XI5/MM1540_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM951 N_NET155_XI5/MM951_d N_NET23_XI5/MM951_g N_VSS_XI5/MM951_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1532 XI5/NET01558 N_NET24_XI5/MM1532_g N_VSS_XI5/MM1532_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM936 N_NET155_XI5/MM936_d N_NET25_XI5/MM936_g N_VSS_XI5/MM936_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1524 XI5/NET01590 N_NET26_XI5/MM1524_g N_VSS_XI5/MM1524_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM919 N_NET155_XI5/MM919_d N_NET27_XI5/MM919_g N_VSS_XI5/MM919_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1516 XI5/NET01622 N_NET28_XI5/MM1516_g N_VSS_XI5/MM1516_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM904 N_NET155_XI5/MM904_d N_NET29_XI5/MM904_g N_VSS_XI5/MM904_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1508 XI5/NET01654 N_NET30_XI5/MM1508_g N_VSS_XI5/MM1508_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM887 N_NET155_XI5/MM887_d N_NET31_XI5/MM887_g N_VSS_XI5/MM887_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1500 XI5/NET01686 N_NET32_XI5/MM1500_g N_VSS_XI5/MM1500_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM872 N_NET155_XI5/MM872_d N_NET33_XI5/MM872_g N_VSS_XI5/MM872_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1492 XI5/NET01718 N_NET34_XI5/MM1492_g N_VSS_XI5/MM1492_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM855 N_NET155_XI5/MM855_d N_NET35_XI5/MM855_g N_VSS_XI5/MM855_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1484 XI5/NET01750 N_NET36_XI5/MM1484_g N_VSS_XI5/MM1484_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM840 N_NET155_XI5/MM840_d N_NET37_XI5/MM840_g N_VSS_XI5/MM840_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1476 XI5/NET01782 N_NET38_XI5/MM1476_g N_VSS_XI5/MM1476_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM823 N_NET155_XI5/MM823_d N_NET39_XI5/MM823_g N_VSS_XI5/MM823_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1468 XI5/NET01814 N_NET40_XI5/MM1468_g N_VSS_XI5/MM1468_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM808 N_NET155_XI5/MM808_d N_NET41_XI5/MM808_g N_VSS_XI5/MM808_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1460 XI5/NET01846 N_NET42_XI5/MM1460_g N_VSS_XI5/MM1460_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM791 N_NET155_XI5/MM791_d N_NET43_XI5/MM791_g N_VSS_XI5/MM791_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1452 XI5/NET01878 N_NET44_XI5/MM1452_g N_VSS_XI5/MM1452_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM776 N_NET155_XI5/MM776_d N_NET45_XI5/MM776_g N_VSS_XI5/MM776_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1444 XI5/NET01910 N_NET46_XI5/MM1444_g N_VSS_XI5/MM1444_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM759 N_NET155_XI5/MM759_d N_NET47_XI5/MM759_g N_VSS_XI5/MM759_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1436 XI5/NET01942 N_NET48_XI5/MM1436_g N_VSS_XI5/MM1436_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM744 N_NET155_XI5/MM744_d N_NET49_XI5/MM744_g N_VSS_XI5/MM744_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1428 XI5/NET01974 N_NET50_XI5/MM1428_g N_VSS_XI5/MM1428_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM728 N_NET155_XI5/MM728_d N_NET51_XI5/MM728_g N_VSS_XI5/MM728_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1420 XI5/NET02006 N_NET52_XI5/MM1420_g N_VSS_XI5/MM1420_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM711 N_NET155_XI5/MM711_d N_NET53_XI5/MM711_g N_VSS_XI5/MM711_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1412 XI5/NET02038 N_NET54_XI5/MM1412_g N_VSS_XI5/MM1412_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM696 N_NET155_XI5/MM696_d N_NET55_XI5/MM696_g N_VSS_XI5/MM696_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1404 XI5/NET02070 N_NET56_XI5/MM1404_g N_VSS_XI5/MM1404_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM679 N_NET155_XI5/MM679_d N_NET57_XI5/MM679_g N_VSS_XI5/MM679_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1396 XI5/NET02102 N_NET58_XI5/MM1396_g N_VSS_XI5/MM1396_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM664 N_NET155_XI5/MM664_d N_NET59_XI5/MM664_g N_VSS_XI5/MM664_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1388 XI5/NET02134 N_NET60_XI5/MM1388_g N_VSS_XI5/MM1388_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM647 N_NET155_XI5/MM647_d N_NET61_XI5/MM647_g N_VSS_XI5/MM647_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1380 XI5/NET02166 N_NET62_XI5/MM1380_g N_VSS_XI5/MM1380_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM632 N_NET155_XI5/MM632_d N_NET63_XI5/MM632_g N_VSS_XI5/MM632_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1372 XI5/NET02198 N_NET64_XI5/MM1372_g N_VSS_XI5/MM1372_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM615 N_NET155_XI5/MM615_d N_NET65_XI5/MM615_g N_VSS_XI5/MM615_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1364 XI5/NET02230 N_NET66_XI5/MM1364_g N_VSS_XI5/MM1364_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM598 N_NET155_XI5/MM598_d N_NET67_XI5/MM598_g N_VSS_XI5/MM598_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1356 XI5/NET02262 N_NET68_XI5/MM1356_g N_VSS_XI5/MM1356_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM585 N_NET155_XI5/MM585_d N_NET69_XI5/MM585_g N_VSS_XI5/MM585_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1348 XI5/NET02294 N_NET70_XI5/MM1348_g N_VSS_XI5/MM1348_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM539 N_NET155_XI5/MM539_d N_NET71_XI5/MM539_g N_VSS_XI5/MM539_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1068 XI5/NET04518 N_NET72_XI5/MM1068_g N_VSS_XI5/MM1068_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM516 N_NET155_XI5/MM516_d N_NET8_XI5/MM516_g N_VSS_XI5/MM516_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI50/MM0 N_NET0215_XI50/MM0_d N_NET0214_XI50/MM0_g N_VSS_XI50/MM0_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI51/MM0 N_NET0214_XI51/MM0_d N_NET134_XI51/MM0_g N_VSS_XI51/MM0_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI7/MM47 N_NET156_XI7/MM47_d N_NET120_XI7/MM47_g N_XI7/NET29_XI7/MM47_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI5/MM1052 N_NET156_XI5/MM1052_d N_NET10_XI5/MM1052_g N_VSS_XI5/MM1052_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1331 XI5/NET02330 N_NET11_XI5/MM1331_g N_VSS_XI5/MM1331_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1027 N_NET156_XI5/MM1027_d N_NET12_XI5/MM1027_g N_VSS_XI5/MM1027_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1325 XI5/NET02354 N_NET13_XI5/MM1325_g N_VSS_XI5/MM1325_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1020 N_NET156_XI5/MM1020_d N_NET14_XI5/MM1020_g N_VSS_XI5/MM1020_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1317 XI5/NET02386 N_NET15_XI5/MM1317_g N_VSS_XI5/MM1317_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM995 N_NET156_XI5/MM995_d N_NET16_XI5/MM995_g N_VSS_XI5/MM995_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1309 XI5/NET02418 N_NET17_XI5/MM1309_g N_VSS_XI5/MM1309_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM988 N_NET156_XI5/MM988_d N_NET18_XI5/MM988_g N_VSS_XI5/MM988_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1301 XI5/NET02450 N_NET19_XI5/MM1301_g N_VSS_XI5/MM1301_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM963 N_NET156_XI5/MM963_d N_NET20_XI5/MM963_g N_VSS_XI5/MM963_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1293 XI5/NET04270 N_NET21_XI5/MM1293_g N_VSS_XI5/MM1293_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM956 N_NET156_XI5/MM956_d N_NET22_XI5/MM956_g N_VSS_XI5/MM956_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1285 XI5/NET04302 N_NET23_XI5/MM1285_g N_VSS_XI5/MM1285_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM931 N_NET156_XI5/MM931_d N_NET24_XI5/MM931_g N_VSS_XI5/MM931_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1277 XI5/NET03450 N_NET25_XI5/MM1277_g N_VSS_XI5/MM1277_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM924 N_NET156_XI5/MM924_d N_NET26_XI5/MM924_g N_VSS_XI5/MM924_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1268 XI5/NET05390 N_NET27_XI5/MM1268_g N_VSS_XI5/MM1268_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM899 N_NET156_XI5/MM899_d N_NET28_XI5/MM899_g N_VSS_XI5/MM899_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1260 XI5/NET05346 N_NET29_XI5/MM1260_g N_VSS_XI5/MM1260_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM892 N_NET156_XI5/MM892_d N_NET30_XI5/MM892_g N_VSS_XI5/MM892_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1252 XI5/NET05302 N_NET31_XI5/MM1252_g N_VSS_XI5/MM1252_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM867 N_NET156_XI5/MM867_d N_NET32_XI5/MM867_g N_VSS_XI5/MM867_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1244 XI5/NET05270 N_NET33_XI5/MM1244_g N_VSS_XI5/MM1244_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM860 N_NET156_XI5/MM860_d N_NET34_XI5/MM860_g N_VSS_XI5/MM860_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1236 XI5/NET05238 N_NET35_XI5/MM1236_g N_VSS_XI5/MM1236_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM835 N_NET156_XI5/MM835_d N_NET36_XI5/MM835_g N_VSS_XI5/MM835_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1228 XI5/NET05206 N_NET37_XI5/MM1228_g N_VSS_XI5/MM1228_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM828 N_NET156_XI5/MM828_d N_NET38_XI5/MM828_g N_VSS_XI5/MM828_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1220 XI5/NET05166 N_NET39_XI5/MM1220_g N_VSS_XI5/MM1220_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM803 N_NET156_XI5/MM803_d N_NET40_XI5/MM803_g N_VSS_XI5/MM803_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1212 XI5/NET05134 N_NET41_XI5/MM1212_g N_VSS_XI5/MM1212_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM796 N_NET156_XI5/MM796_d N_NET42_XI5/MM796_g N_VSS_XI5/MM796_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1204 XI5/NET05098 N_NET43_XI5/MM1204_g N_VSS_XI5/MM1204_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM771 N_NET156_XI5/MM771_d N_NET44_XI5/MM771_g N_VSS_XI5/MM771_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1196 XI5/NET05066 N_NET45_XI5/MM1196_g N_VSS_XI5/MM1196_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM764 N_NET156_XI5/MM764_d N_NET46_XI5/MM764_g N_VSS_XI5/MM764_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1188 XI5/NET05034 N_NET47_XI5/MM1188_g N_VSS_XI5/MM1188_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM739 N_NET156_XI5/MM739_d N_NET48_XI5/MM739_g N_VSS_XI5/MM739_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1180 XI5/NET05002 N_NET49_XI5/MM1180_g N_VSS_XI5/MM1180_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM723 N_NET156_XI5/MM723_d N_NET50_XI5/MM723_g N_VSS_XI5/MM723_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1172 XI5/NET04970 N_NET51_XI5/MM1172_g N_VSS_XI5/MM1172_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM716 N_NET156_XI5/MM716_d N_NET52_XI5/MM716_g N_VSS_XI5/MM716_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1164 XI5/NET04938 N_NET53_XI5/MM1164_g N_VSS_XI5/MM1164_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM691 N_NET156_XI5/MM691_d N_NET54_XI5/MM691_g N_VSS_XI5/MM691_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1156 XI5/NET04898 N_NET55_XI5/MM1156_g N_VSS_XI5/MM1156_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM684 N_NET156_XI5/MM684_d N_NET56_XI5/MM684_g N_VSS_XI5/MM684_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1148 XI5/NET04866 N_NET57_XI5/MM1148_g N_VSS_XI5/MM1148_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM659 N_NET156_XI5/MM659_d N_NET58_XI5/MM659_g N_VSS_XI5/MM659_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1140 XI5/NET04834 N_NET59_XI5/MM1140_g N_VSS_XI5/MM1140_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM652 N_NET156_XI5/MM652_d N_NET60_XI5/MM652_g N_VSS_XI5/MM652_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1132 XI5/NET04802 N_NET61_XI5/MM1132_g N_VSS_XI5/MM1132_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM627 N_NET156_XI5/MM627_d N_NET62_XI5/MM627_g N_VSS_XI5/MM627_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1124 XI5/NET04750 N_NET63_XI5/MM1124_g N_VSS_XI5/MM1124_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM620 N_NET156_XI5/MM620_d N_NET64_XI5/MM620_g N_VSS_XI5/MM620_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1107 XI5/NET04710 N_NET65_XI5/MM1107_g N_VSS_XI5/MM1107_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM603 N_NET156_XI5/MM603_d N_NET66_XI5/MM603_g N_VSS_XI5/MM603_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1091 XI5/NET04634 N_NET67_XI5/MM1091_g N_VSS_XI5/MM1091_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM580 N_NET156_XI5/MM580_d N_NET68_XI5/MM580_g N_VSS_XI5/MM580_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1083 XI5/NET04602 N_NET69_XI5/MM1083_g N_VSS_XI5/MM1083_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM537 N_NET156_XI5/MM537_d N_NET70_XI5/MM537_g N_VSS_XI5/MM537_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1075 XI5/NET04558 N_NET71_XI5/MM1075_g N_VSS_XI5/MM1075_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM522 N_NET156_XI5/MM522_d N_NET72_XI5/MM522_g N_VSS_XI5/MM522_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1059 XI5/NET04370 N_NET8_XI5/MM1059_g N_VSS_XI5/MM1059_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM46 N_NET157_XI7/MM46_d N_XI7/NET48_XI7/MM46_g N_XI7/NET29_XI7/MM46_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI5/MM1589 XI5/NET01330 N_NET10_XI5/MM1589_g N_VSS_XI5/MM1589_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1048 N_NET157_XI5/MM1048_d N_NET11_XI5/MM1048_g N_VSS_XI5/MM1048_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1581 XI5/NET01362 N_NET12_XI5/MM1581_g N_VSS_XI5/MM1581_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1031 N_NET157_XI5/MM1031_d N_NET13_XI5/MM1031_g N_VSS_XI5/MM1031_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1573 XI5/NET01394 N_NET14_XI5/MM1573_g N_VSS_XI5/MM1573_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1016 N_NET157_XI5/MM1016_d N_NET15_XI5/MM1016_g N_VSS_XI5/MM1016_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1565 XI5/NET01426 N_NET16_XI5/MM1565_g N_VSS_XI5/MM1565_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM999 N_NET157_XI5/MM999_d N_NET17_XI5/MM999_g N_VSS_XI5/MM999_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1557 XI5/NET01458 N_NET18_XI5/MM1557_g N_VSS_XI5/MM1557_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM984 N_NET157_XI5/MM984_d N_NET19_XI5/MM984_g N_VSS_XI5/MM984_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1549 XI5/NET01490 N_NET20_XI5/MM1549_g N_VSS_XI5/MM1549_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM967 N_NET157_XI5/MM967_d N_NET21_XI5/MM967_g N_VSS_XI5/MM967_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1541 XI5/NET01522 N_NET22_XI5/MM1541_g N_VSS_XI5/MM1541_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM952 N_NET157_XI5/MM952_d N_NET23_XI5/MM952_g N_VSS_XI5/MM952_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1533 XI5/NET01554 N_NET24_XI5/MM1533_g N_VSS_XI5/MM1533_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM935 N_NET157_XI5/MM935_d N_NET25_XI5/MM935_g N_VSS_XI5/MM935_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1525 XI5/NET01586 N_NET26_XI5/MM1525_g N_VSS_XI5/MM1525_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM920 N_NET157_XI5/MM920_d N_NET27_XI5/MM920_g N_VSS_XI5/MM920_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1517 XI5/NET01618 N_NET28_XI5/MM1517_g N_VSS_XI5/MM1517_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM903 N_NET157_XI5/MM903_d N_NET29_XI5/MM903_g N_VSS_XI5/MM903_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1509 XI5/NET01650 N_NET30_XI5/MM1509_g N_VSS_XI5/MM1509_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM888 N_NET157_XI5/MM888_d N_NET31_XI5/MM888_g N_VSS_XI5/MM888_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1501 XI5/NET01682 N_NET32_XI5/MM1501_g N_VSS_XI5/MM1501_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM871 N_NET157_XI5/MM871_d N_NET33_XI5/MM871_g N_VSS_XI5/MM871_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1493 XI5/NET01714 N_NET34_XI5/MM1493_g N_VSS_XI5/MM1493_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM856 N_NET157_XI5/MM856_d N_NET35_XI5/MM856_g N_VSS_XI5/MM856_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1485 XI5/NET01746 N_NET36_XI5/MM1485_g N_VSS_XI5/MM1485_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM839 N_NET157_XI5/MM839_d N_NET37_XI5/MM839_g N_VSS_XI5/MM839_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1477 XI5/NET01778 N_NET38_XI5/MM1477_g N_VSS_XI5/MM1477_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM824 N_NET157_XI5/MM824_d N_NET39_XI5/MM824_g N_VSS_XI5/MM824_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1469 XI5/NET01810 N_NET40_XI5/MM1469_g N_VSS_XI5/MM1469_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM807 N_NET157_XI5/MM807_d N_NET41_XI5/MM807_g N_VSS_XI5/MM807_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1461 XI5/NET01842 N_NET42_XI5/MM1461_g N_VSS_XI5/MM1461_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM792 N_NET157_XI5/MM792_d N_NET43_XI5/MM792_g N_VSS_XI5/MM792_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1453 XI5/NET01874 N_NET44_XI5/MM1453_g N_VSS_XI5/MM1453_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM775 N_NET157_XI5/MM775_d N_NET45_XI5/MM775_g N_VSS_XI5/MM775_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1445 XI5/NET01906 N_NET46_XI5/MM1445_g N_VSS_XI5/MM1445_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM760 N_NET157_XI5/MM760_d N_NET47_XI5/MM760_g N_VSS_XI5/MM760_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1437 XI5/NET01938 N_NET48_XI5/MM1437_g N_VSS_XI5/MM1437_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM743 N_NET157_XI5/MM743_d N_NET49_XI5/MM743_g N_VSS_XI5/MM743_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1429 XI5/NET01970 N_NET50_XI5/MM1429_g N_VSS_XI5/MM1429_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM727 N_NET157_XI5/MM727_d N_NET51_XI5/MM727_g N_VSS_XI5/MM727_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1421 XI5/NET02002 N_NET52_XI5/MM1421_g N_VSS_XI5/MM1421_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM712 N_NET157_XI5/MM712_d N_NET53_XI5/MM712_g N_VSS_XI5/MM712_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1413 XI5/NET02034 N_NET54_XI5/MM1413_g N_VSS_XI5/MM1413_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM695 N_NET157_XI5/MM695_d N_NET55_XI5/MM695_g N_VSS_XI5/MM695_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1405 XI5/NET02066 N_NET56_XI5/MM1405_g N_VSS_XI5/MM1405_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM680 N_NET157_XI5/MM680_d N_NET57_XI5/MM680_g N_VSS_XI5/MM680_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1397 XI5/NET02098 N_NET58_XI5/MM1397_g N_VSS_XI5/MM1397_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM663 N_NET157_XI5/MM663_d N_NET59_XI5/MM663_g N_VSS_XI5/MM663_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1389 XI5/NET02130 N_NET60_XI5/MM1389_g N_VSS_XI5/MM1389_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM648 N_NET157_XI5/MM648_d N_NET61_XI5/MM648_g N_VSS_XI5/MM648_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1381 XI5/NET02162 N_NET62_XI5/MM1381_g N_VSS_XI5/MM1381_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM631 N_NET157_XI5/MM631_d N_NET63_XI5/MM631_g N_VSS_XI5/MM631_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1373 XI5/NET02194 N_NET64_XI5/MM1373_g N_VSS_XI5/MM1373_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM616 N_NET157_XI5/MM616_d N_NET65_XI5/MM616_g N_VSS_XI5/MM616_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1365 XI5/NET02226 N_NET66_XI5/MM1365_g N_VSS_XI5/MM1365_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM599 N_NET157_XI5/MM599_d N_NET67_XI5/MM599_g N_VSS_XI5/MM599_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1357 XI5/NET02258 N_NET68_XI5/MM1357_g N_VSS_XI5/MM1357_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM584 N_NET157_XI5/MM584_d N_NET69_XI5/MM584_g N_VSS_XI5/MM584_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1350 XI5/NET02286 N_NET70_XI5/MM1350_g N_VSS_XI5/MM1350_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM538 N_NET157_XI5/MM538_d N_NET71_XI5/MM538_g N_VSS_XI5/MM538_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1067 XI5/NET04514 N_NET72_XI5/MM1067_g N_VSS_XI5/MM1067_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM518 N_NET157_XI5/MM518_d N_NET8_XI5/MM518_g N_VSS_XI5/MM518_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM38 N_XI7/NET29_XI7/MM38_d N_NET125_XI7/MM38_g N_XI7/NET57_XI7/MM38_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI9/MM1 N_NET134_XI9/MM1_d N_NET0181_XI9/MM1_g N_XI9/NET40_XI9/MM1_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=1e-06 AD=5e-13 AS=1.5e-13 PD=2e-06
+ PS=3e-07
mXI9/MM0 N_XI9/NET40_XI9/MM0_d N_VREF_XI9/MM0_g N_XI9/NET43_XI9/MM0_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=1e-06 AD=1.5e-13 AS=2.7e-13 PD=3e-07
+ PS=5.4e-07
mXI9/MM4 N_XI9/NET43_XI9/MM4_d N_NET82_XI9/MM4_g N_VSS_XI9/MM4_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=1e-06 AD=2.7e-13 AS=2.55e-13
+ PD=5.4e-07 PS=5.1e-07
mXI9/MM4@2 N_XI9/NET43_XI9/MM4@2_d N_NET82_XI9/MM4@2_g N_VSS_XI9/MM4@2_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=1e-06 AD=2.7e-13 AS=2.55e-13
+ PD=5.4e-07 PS=5.1e-07
mXI9/MM3 N_XI9/NET28_XI9/MM3_d N_NET165_XI9/MM3_g N_XI9/NET43_XI9/MM3_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=1e-06 AD=1.725e-13 AS=2.7e-13
+ PD=3.45e-07 PS=5.4e-07
mXI9/MM2 N_NET0181_XI9/MM2_d N_NET134_XI9/MM2_g N_XI9/NET28_XI9/MM2_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=1.725e-13
+ PD=1.98e-06 PS=3.45e-07
mXI7/MM39 N_XI7/NET33_XI7/MM39_d N_XI7/NET68_XI7/MM39_g N_XI7/NET57_XI7/MM39_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI7/MM44 N_NET150_XI7/MM44_d N_NET120_XI7/MM44_g N_XI7/NET33_XI7/MM44_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI5/MM1050 N_NET150_XI5/MM1050_d N_NET10_XI5/MM1050_g N_VSS_XI5/MM1050_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1335 XI5/NET02314 N_NET11_XI5/MM1335_g N_VSS_XI5/MM1335_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1029 N_NET150_XI5/MM1029_d N_NET12_XI5/MM1029_g N_VSS_XI5/MM1029_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1326 XI5/NET02350 N_NET13_XI5/MM1326_g N_VSS_XI5/MM1326_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1018 N_NET150_XI5/MM1018_d N_NET14_XI5/MM1018_g N_VSS_XI5/MM1018_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1318 XI5/NET02382 N_NET15_XI5/MM1318_g N_VSS_XI5/MM1318_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM997 N_NET150_XI5/MM997_d N_NET16_XI5/MM997_g N_VSS_XI5/MM997_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1310 XI5/NET02414 N_NET17_XI5/MM1310_g N_VSS_XI5/MM1310_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM986 N_NET150_XI5/MM986_d N_NET18_XI5/MM986_g N_VSS_XI5/MM986_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1302 XI5/NET02446 N_NET19_XI5/MM1302_g N_VSS_XI5/MM1302_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM965 N_NET150_XI5/MM965_d N_NET20_XI5/MM965_g N_VSS_XI5/MM965_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1294 XI5/NET04266 N_NET21_XI5/MM1294_g N_VSS_XI5/MM1294_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM954 N_NET150_XI5/MM954_d N_NET22_XI5/MM954_g N_VSS_XI5/MM954_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1286 XI5/NET04298 N_NET23_XI5/MM1286_g N_VSS_XI5/MM1286_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM933 N_NET150_XI5/MM933_d N_NET24_XI5/MM933_g N_VSS_XI5/MM933_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1278 XI5/NET03446 N_NET25_XI5/MM1278_g N_VSS_XI5/MM1278_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM922 N_NET150_XI5/MM922_d N_NET26_XI5/MM922_g N_VSS_XI5/MM922_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1267 XI5/NET05386 N_NET27_XI5/MM1267_g N_VSS_XI5/MM1267_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM901 N_NET150_XI5/MM901_d N_NET28_XI5/MM901_g N_VSS_XI5/MM901_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1259 XI5/NET05342 N_NET29_XI5/MM1259_g N_VSS_XI5/MM1259_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM890 N_NET150_XI5/MM890_d N_NET30_XI5/MM890_g N_VSS_XI5/MM890_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1251 XI5/NET05298 N_NET31_XI5/MM1251_g N_VSS_XI5/MM1251_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM869 N_NET150_XI5/MM869_d N_NET32_XI5/MM869_g N_VSS_XI5/MM869_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1243 XI5/NET05266 N_NET33_XI5/MM1243_g N_VSS_XI5/MM1243_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM858 N_NET150_XI5/MM858_d N_NET34_XI5/MM858_g N_VSS_XI5/MM858_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1235 XI5/NET05234 N_NET35_XI5/MM1235_g N_VSS_XI5/MM1235_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM837 N_NET150_XI5/MM837_d N_NET36_XI5/MM837_g N_VSS_XI5/MM837_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1227 XI5/NET05202 N_NET37_XI5/MM1227_g N_VSS_XI5/MM1227_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM826 N_NET150_XI5/MM826_d N_NET38_XI5/MM826_g N_VSS_XI5/MM826_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1219 XI5/NET05162 N_NET39_XI5/MM1219_g N_VSS_XI5/MM1219_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM805 N_NET150_XI5/MM805_d N_NET40_XI5/MM805_g N_VSS_XI5/MM805_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1211 XI5/NET05130 N_NET41_XI5/MM1211_g N_VSS_XI5/MM1211_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM794 N_NET150_XI5/MM794_d N_NET42_XI5/MM794_g N_VSS_XI5/MM794_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1203 XI5/NET05094 N_NET43_XI5/MM1203_g N_VSS_XI5/MM1203_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM773 N_NET150_XI5/MM773_d N_NET44_XI5/MM773_g N_VSS_XI5/MM773_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1195 XI5/NET05062 N_NET45_XI5/MM1195_g N_VSS_XI5/MM1195_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM762 N_NET150_XI5/MM762_d N_NET46_XI5/MM762_g N_VSS_XI5/MM762_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1187 XI5/NET05030 N_NET47_XI5/MM1187_g N_VSS_XI5/MM1187_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM741 N_NET150_XI5/MM741_d N_NET48_XI5/MM741_g N_VSS_XI5/MM741_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1179 XI5/NET04998 N_NET49_XI5/MM1179_g N_VSS_XI5/MM1179_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM725 N_NET150_XI5/MM725_d N_NET50_XI5/MM725_g N_VSS_XI5/MM725_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1171 XI5/NET04966 N_NET51_XI5/MM1171_g N_VSS_XI5/MM1171_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM714 N_NET150_XI5/MM714_d N_NET52_XI5/MM714_g N_VSS_XI5/MM714_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1163 XI5/NET04934 N_NET53_XI5/MM1163_g N_VSS_XI5/MM1163_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM693 N_NET150_XI5/MM693_d N_NET54_XI5/MM693_g N_VSS_XI5/MM693_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1155 XI5/NET04894 N_NET55_XI5/MM1155_g N_VSS_XI5/MM1155_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM682 N_NET150_XI5/MM682_d N_NET56_XI5/MM682_g N_VSS_XI5/MM682_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1147 XI5/NET04862 N_NET57_XI5/MM1147_g N_VSS_XI5/MM1147_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM661 N_NET150_XI5/MM661_d N_NET58_XI5/MM661_g N_VSS_XI5/MM661_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1139 XI5/NET04830 N_NET59_XI5/MM1139_g N_VSS_XI5/MM1139_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM650 N_NET150_XI5/MM650_d N_NET60_XI5/MM650_g N_VSS_XI5/MM650_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1131 XI5/NET04798 N_NET61_XI5/MM1131_g N_VSS_XI5/MM1131_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM629 N_NET150_XI5/MM629_d N_NET62_XI5/MM629_g N_VSS_XI5/MM629_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1123 XI5/NET04746 N_NET63_XI5/MM1123_g N_VSS_XI5/MM1123_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM618 N_NET150_XI5/MM618_d N_NET64_XI5/MM618_g N_VSS_XI5/MM618_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1106 XI5/NET04706 N_NET65_XI5/MM1106_g N_VSS_XI5/MM1106_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM601 N_NET150_XI5/MM601_d N_NET66_XI5/MM601_g N_VSS_XI5/MM601_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1090 XI5/NET04630 N_NET67_XI5/MM1090_g N_VSS_XI5/MM1090_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM582 N_NET150_XI5/MM582_d N_NET68_XI5/MM582_g N_VSS_XI5/MM582_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1082 XI5/NET04598 N_NET69_XI5/MM1082_g N_VSS_XI5/MM1082_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM532 N_NET150_XI5/MM532_d N_NET70_XI5/MM532_g N_VSS_XI5/MM532_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1074 XI5/NET04554 N_NET71_XI5/MM1074_g N_VSS_XI5/MM1074_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM527 N_NET150_XI5/MM527_d N_NET72_XI5/MM527_g N_VSS_XI5/MM527_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1058 XI5/NET04322 N_NET8_XI5/MM1058_g N_VSS_XI5/MM1058_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM45 N_NET158_XI7/MM45_d N_XI7/NET48_XI7/MM45_g N_XI7/NET33_XI7/MM45_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI5/MM1590 XI5/NET01326 N_NET10_XI5/MM1590_g N_VSS_XI5/MM1590_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1043 N_NET158_XI5/MM1043_d N_NET11_XI5/MM1043_g N_VSS_XI5/MM1043_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1582 XI5/NET01358 N_NET12_XI5/MM1582_g N_VSS_XI5/MM1582_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1036 N_NET158_XI5/MM1036_d N_NET13_XI5/MM1036_g N_VSS_XI5/MM1036_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1574 XI5/NET01390 N_NET14_XI5/MM1574_g N_VSS_XI5/MM1574_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1011 N_NET158_XI5/MM1011_d N_NET15_XI5/MM1011_g N_VSS_XI5/MM1011_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1566 XI5/NET01422 N_NET16_XI5/MM1566_g N_VSS_XI5/MM1566_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1004 N_NET158_XI5/MM1004_d N_NET17_XI5/MM1004_g N_VSS_XI5/MM1004_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1558 XI5/NET01454 N_NET18_XI5/MM1558_g N_VSS_XI5/MM1558_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM979 N_NET158_XI5/MM979_d N_NET19_XI5/MM979_g N_VSS_XI5/MM979_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1550 XI5/NET01486 N_NET20_XI5/MM1550_g N_VSS_XI5/MM1550_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM972 N_NET158_XI5/MM972_d N_NET21_XI5/MM972_g N_VSS_XI5/MM972_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1542 XI5/NET01518 N_NET22_XI5/MM1542_g N_VSS_XI5/MM1542_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM947 N_NET158_XI5/MM947_d N_NET23_XI5/MM947_g N_VSS_XI5/MM947_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1534 XI5/NET01550 N_NET24_XI5/MM1534_g N_VSS_XI5/MM1534_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM940 N_NET158_XI5/MM940_d N_NET25_XI5/MM940_g N_VSS_XI5/MM940_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1526 XI5/NET01582 N_NET26_XI5/MM1526_g N_VSS_XI5/MM1526_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM915 N_NET158_XI5/MM915_d N_NET27_XI5/MM915_g N_VSS_XI5/MM915_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1518 XI5/NET01614 N_NET28_XI5/MM1518_g N_VSS_XI5/MM1518_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM908 N_NET158_XI5/MM908_d N_NET29_XI5/MM908_g N_VSS_XI5/MM908_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1510 XI5/NET01646 N_NET30_XI5/MM1510_g N_VSS_XI5/MM1510_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM883 N_NET158_XI5/MM883_d N_NET31_XI5/MM883_g N_VSS_XI5/MM883_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1502 XI5/NET01678 N_NET32_XI5/MM1502_g N_VSS_XI5/MM1502_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM876 N_NET158_XI5/MM876_d N_NET33_XI5/MM876_g N_VSS_XI5/MM876_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1494 XI5/NET01710 N_NET34_XI5/MM1494_g N_VSS_XI5/MM1494_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM851 N_NET158_XI5/MM851_d N_NET35_XI5/MM851_g N_VSS_XI5/MM851_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1486 XI5/NET01742 N_NET36_XI5/MM1486_g N_VSS_XI5/MM1486_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM844 N_NET158_XI5/MM844_d N_NET37_XI5/MM844_g N_VSS_XI5/MM844_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1478 XI5/NET01774 N_NET38_XI5/MM1478_g N_VSS_XI5/MM1478_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM819 N_NET158_XI5/MM819_d N_NET39_XI5/MM819_g N_VSS_XI5/MM819_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1470 XI5/NET01806 N_NET40_XI5/MM1470_g N_VSS_XI5/MM1470_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM812 N_NET158_XI5/MM812_d N_NET41_XI5/MM812_g N_VSS_XI5/MM812_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1462 XI5/NET01838 N_NET42_XI5/MM1462_g N_VSS_XI5/MM1462_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM787 N_NET158_XI5/MM787_d N_NET43_XI5/MM787_g N_VSS_XI5/MM787_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1454 XI5/NET01870 N_NET44_XI5/MM1454_g N_VSS_XI5/MM1454_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM780 N_NET158_XI5/MM780_d N_NET45_XI5/MM780_g N_VSS_XI5/MM780_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1446 XI5/NET01902 N_NET46_XI5/MM1446_g N_VSS_XI5/MM1446_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM755 N_NET158_XI5/MM755_d N_NET47_XI5/MM755_g N_VSS_XI5/MM755_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1438 XI5/NET01934 N_NET48_XI5/MM1438_g N_VSS_XI5/MM1438_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM748 N_NET158_XI5/MM748_d N_NET49_XI5/MM748_g N_VSS_XI5/MM748_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1430 XI5/NET01966 N_NET50_XI5/MM1430_g N_VSS_XI5/MM1430_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM732 N_NET158_XI5/MM732_d N_NET51_XI5/MM732_g N_VSS_XI5/MM732_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1422 XI5/NET01998 N_NET52_XI5/MM1422_g N_VSS_XI5/MM1422_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM707 N_NET158_XI5/MM707_d N_NET53_XI5/MM707_g N_VSS_XI5/MM707_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1414 XI5/NET02030 N_NET54_XI5/MM1414_g N_VSS_XI5/MM1414_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM700 N_NET158_XI5/MM700_d N_NET55_XI5/MM700_g N_VSS_XI5/MM700_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1406 XI5/NET02062 N_NET56_XI5/MM1406_g N_VSS_XI5/MM1406_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM675 N_NET158_XI5/MM675_d N_NET57_XI5/MM675_g N_VSS_XI5/MM675_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1398 XI5/NET02094 N_NET58_XI5/MM1398_g N_VSS_XI5/MM1398_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM668 N_NET158_XI5/MM668_d N_NET59_XI5/MM668_g N_VSS_XI5/MM668_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1390 XI5/NET02126 N_NET60_XI5/MM1390_g N_VSS_XI5/MM1390_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM643 N_NET158_XI5/MM643_d N_NET61_XI5/MM643_g N_VSS_XI5/MM643_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1382 XI5/NET02158 N_NET62_XI5/MM1382_g N_VSS_XI5/MM1382_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM636 N_NET158_XI5/MM636_d N_NET63_XI5/MM636_g N_VSS_XI5/MM636_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1374 XI5/NET02190 N_NET64_XI5/MM1374_g N_VSS_XI5/MM1374_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM611 N_NET158_XI5/MM611_d N_NET65_XI5/MM611_g N_VSS_XI5/MM611_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1366 XI5/NET02222 N_NET66_XI5/MM1366_g N_VSS_XI5/MM1366_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM594 N_NET158_XI5/MM594_d N_NET67_XI5/MM594_g N_VSS_XI5/MM594_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1358 XI5/NET02254 N_NET68_XI5/MM1358_g N_VSS_XI5/MM1358_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM589 N_NET158_XI5/MM589_d N_NET69_XI5/MM589_g N_VSS_XI5/MM589_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1345 XI5/NET02306 N_NET70_XI5/MM1345_g N_VSS_XI5/MM1345_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM543 N_NET158_XI5/MM543_d N_NET71_XI5/MM543_g N_VSS_XI5/MM543_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1066 XI5/NET04510 N_NET72_XI5/MM1066_g N_VSS_XI5/MM1066_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM519 N_NET158_XI5/MM519_d N_NET8_XI5/MM519_g N_VSS_XI5/MM519_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM35 N_XI7/NET57_XI7/MM35_d N_NET85_XI7/MM35_g N_NET165_XI7/MM35_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI7/MM34 N_XI7/NET69_XI7/MM34_d N_XI7/NET76_XI7/MM34_g N_NET165_XI7/MM34_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI7/MM43 N_NET159_XI7/MM43_d N_NET120_XI7/MM43_g N_XI7/NET45_XI7/MM43_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI5/MM1054 N_NET159_XI5/MM1054_d N_NET10_XI5/MM1054_g N_VSS_XI5/MM1054_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1334 XI5/NET02318 N_NET11_XI5/MM1334_g N_VSS_XI5/MM1334_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1025 N_NET159_XI5/MM1025_d N_NET12_XI5/MM1025_g N_VSS_XI5/MM1025_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1327 XI5/NET02346 N_NET13_XI5/MM1327_g N_VSS_XI5/MM1327_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1022 N_NET159_XI5/MM1022_d N_NET14_XI5/MM1022_g N_VSS_XI5/MM1022_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1319 XI5/NET02378 N_NET15_XI5/MM1319_g N_VSS_XI5/MM1319_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM993 N_NET159_XI5/MM993_d N_NET16_XI5/MM993_g N_VSS_XI5/MM993_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1311 XI5/NET02410 N_NET17_XI5/MM1311_g N_VSS_XI5/MM1311_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM990 N_NET159_XI5/MM990_d N_NET18_XI5/MM990_g N_VSS_XI5/MM990_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1303 XI5/NET02442 N_NET19_XI5/MM1303_g N_VSS_XI5/MM1303_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM961 N_NET159_XI5/MM961_d N_NET20_XI5/MM961_g N_VSS_XI5/MM961_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1295 XI5/NET04262 N_NET21_XI5/MM1295_g N_VSS_XI5/MM1295_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM958 N_NET159_XI5/MM958_d N_NET22_XI5/MM958_g N_VSS_XI5/MM958_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1287 XI5/NET04294 N_NET23_XI5/MM1287_g N_VSS_XI5/MM1287_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM929 N_NET159_XI5/MM929_d N_NET24_XI5/MM929_g N_VSS_XI5/MM929_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1279 XI5/NET03442 N_NET25_XI5/MM1279_g N_VSS_XI5/MM1279_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM926 N_NET159_XI5/MM926_d N_NET26_XI5/MM926_g N_VSS_XI5/MM926_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1266 XI5/NET05382 N_NET27_XI5/MM1266_g N_VSS_XI5/MM1266_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM897 N_NET159_XI5/MM897_d N_NET28_XI5/MM897_g N_VSS_XI5/MM897_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1258 XI5/NET05338 N_NET29_XI5/MM1258_g N_VSS_XI5/MM1258_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM894 N_NET159_XI5/MM894_d N_NET30_XI5/MM894_g N_VSS_XI5/MM894_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1250 XI5/NET05294 N_NET31_XI5/MM1250_g N_VSS_XI5/MM1250_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM865 N_NET159_XI5/MM865_d N_NET32_XI5/MM865_g N_VSS_XI5/MM865_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1242 XI5/NET05262 N_NET33_XI5/MM1242_g N_VSS_XI5/MM1242_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM862 N_NET159_XI5/MM862_d N_NET34_XI5/MM862_g N_VSS_XI5/MM862_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1234 XI5/NET05230 N_NET35_XI5/MM1234_g N_VSS_XI5/MM1234_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM833 N_NET159_XI5/MM833_d N_NET36_XI5/MM833_g N_VSS_XI5/MM833_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1226 XI5/NET05198 N_NET37_XI5/MM1226_g N_VSS_XI5/MM1226_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM830 N_NET159_XI5/MM830_d N_NET38_XI5/MM830_g N_VSS_XI5/MM830_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1218 XI5/NET05158 N_NET39_XI5/MM1218_g N_VSS_XI5/MM1218_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM801 N_NET159_XI5/MM801_d N_NET40_XI5/MM801_g N_VSS_XI5/MM801_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1210 XI5/NET05126 N_NET41_XI5/MM1210_g N_VSS_XI5/MM1210_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM798 N_NET159_XI5/MM798_d N_NET42_XI5/MM798_g N_VSS_XI5/MM798_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1202 XI5/NET05090 N_NET43_XI5/MM1202_g N_VSS_XI5/MM1202_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM769 N_NET159_XI5/MM769_d N_NET44_XI5/MM769_g N_VSS_XI5/MM769_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1194 XI5/NET05058 N_NET45_XI5/MM1194_g N_VSS_XI5/MM1194_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM766 N_NET159_XI5/MM766_d N_NET46_XI5/MM766_g N_VSS_XI5/MM766_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1186 XI5/NET05026 N_NET47_XI5/MM1186_g N_VSS_XI5/MM1186_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM737 N_NET159_XI5/MM737_d N_NET48_XI5/MM737_g N_VSS_XI5/MM737_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1178 XI5/NET04994 N_NET49_XI5/MM1178_g N_VSS_XI5/MM1178_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM721 N_NET159_XI5/MM721_d N_NET50_XI5/MM721_g N_VSS_XI5/MM721_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1170 XI5/NET04962 N_NET51_XI5/MM1170_g N_VSS_XI5/MM1170_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM718 N_NET159_XI5/MM718_d N_NET52_XI5/MM718_g N_VSS_XI5/MM718_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1162 XI5/NET04930 N_NET53_XI5/MM1162_g N_VSS_XI5/MM1162_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM689 N_NET159_XI5/MM689_d N_NET54_XI5/MM689_g N_VSS_XI5/MM689_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1154 XI5/NET04890 N_NET55_XI5/MM1154_g N_VSS_XI5/MM1154_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM686 N_NET159_XI5/MM686_d N_NET56_XI5/MM686_g N_VSS_XI5/MM686_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1146 XI5/NET04858 N_NET57_XI5/MM1146_g N_VSS_XI5/MM1146_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM657 N_NET159_XI5/MM657_d N_NET58_XI5/MM657_g N_VSS_XI5/MM657_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1138 XI5/NET04826 N_NET59_XI5/MM1138_g N_VSS_XI5/MM1138_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM654 N_NET159_XI5/MM654_d N_NET60_XI5/MM654_g N_VSS_XI5/MM654_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1130 XI5/NET04794 N_NET61_XI5/MM1130_g N_VSS_XI5/MM1130_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM625 N_NET159_XI5/MM625_d N_NET62_XI5/MM625_g N_VSS_XI5/MM625_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1121 XI5/NET04742 N_NET63_XI5/MM1121_g N_VSS_XI5/MM1121_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM622 N_NET159_XI5/MM622_d N_NET64_XI5/MM622_g N_VSS_XI5/MM622_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1104 XI5/NET04694 N_NET65_XI5/MM1104_g N_VSS_XI5/MM1104_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM606 N_NET159_XI5/MM606_d N_NET66_XI5/MM606_g N_VSS_XI5/MM606_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1089 XI5/NET04626 N_NET67_XI5/MM1089_g N_VSS_XI5/MM1089_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM577 N_NET159_XI5/MM577_d N_NET68_XI5/MM577_g N_VSS_XI5/MM577_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1081 XI5/NET04594 N_NET69_XI5/MM1081_g N_VSS_XI5/MM1081_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM534 N_NET159_XI5/MM534_d N_NET70_XI5/MM534_g N_VSS_XI5/MM534_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1073 XI5/NET04550 N_NET71_XI5/MM1073_g N_VSS_XI5/MM1073_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM525 N_NET159_XI5/MM525_d N_NET72_XI5/MM525_g N_VSS_XI5/MM525_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1057 XI5/NET03002 N_NET8_XI5/MM1057_g N_VSS_XI5/MM1057_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM42 N_NET160_XI7/MM42_d N_XI7/NET48_XI7/MM42_g N_XI7/NET45_XI7/MM42_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI5/MM1591 XI5/NET01322 N_NET10_XI5/MM1591_g N_VSS_XI5/MM1591_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1045 N_NET160_XI5/MM1045_d N_NET11_XI5/MM1045_g N_VSS_XI5/MM1045_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1583 XI5/NET01354 N_NET12_XI5/MM1583_g N_VSS_XI5/MM1583_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1034 N_NET160_XI5/MM1034_d N_NET13_XI5/MM1034_g N_VSS_XI5/MM1034_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1575 XI5/NET01386 N_NET14_XI5/MM1575_g N_VSS_XI5/MM1575_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1013 N_NET160_XI5/MM1013_d N_NET15_XI5/MM1013_g N_VSS_XI5/MM1013_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1567 XI5/NET01418 N_NET16_XI5/MM1567_g N_VSS_XI5/MM1567_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1002 N_NET160_XI5/MM1002_d N_NET17_XI5/MM1002_g N_VSS_XI5/MM1002_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1559 XI5/NET01450 N_NET18_XI5/MM1559_g N_VSS_XI5/MM1559_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM981 N_NET160_XI5/MM981_d N_NET19_XI5/MM981_g N_VSS_XI5/MM981_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1551 XI5/NET01482 N_NET20_XI5/MM1551_g N_VSS_XI5/MM1551_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM970 N_NET160_XI5/MM970_d N_NET21_XI5/MM970_g N_VSS_XI5/MM970_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1543 XI5/NET01514 N_NET22_XI5/MM1543_g N_VSS_XI5/MM1543_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM949 N_NET160_XI5/MM949_d N_NET23_XI5/MM949_g N_VSS_XI5/MM949_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1535 XI5/NET01546 N_NET24_XI5/MM1535_g N_VSS_XI5/MM1535_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM938 N_NET160_XI5/MM938_d N_NET25_XI5/MM938_g N_VSS_XI5/MM938_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1527 XI5/NET01578 N_NET26_XI5/MM1527_g N_VSS_XI5/MM1527_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM917 N_NET160_XI5/MM917_d N_NET27_XI5/MM917_g N_VSS_XI5/MM917_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1519 XI5/NET01610 N_NET28_XI5/MM1519_g N_VSS_XI5/MM1519_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM906 N_NET160_XI5/MM906_d N_NET29_XI5/MM906_g N_VSS_XI5/MM906_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1511 XI5/NET01642 N_NET30_XI5/MM1511_g N_VSS_XI5/MM1511_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM885 N_NET160_XI5/MM885_d N_NET31_XI5/MM885_g N_VSS_XI5/MM885_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1503 XI5/NET01674 N_NET32_XI5/MM1503_g N_VSS_XI5/MM1503_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM874 N_NET160_XI5/MM874_d N_NET33_XI5/MM874_g N_VSS_XI5/MM874_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1495 XI5/NET01706 N_NET34_XI5/MM1495_g N_VSS_XI5/MM1495_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM853 N_NET160_XI5/MM853_d N_NET35_XI5/MM853_g N_VSS_XI5/MM853_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1487 XI5/NET01738 N_NET36_XI5/MM1487_g N_VSS_XI5/MM1487_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM842 N_NET160_XI5/MM842_d N_NET37_XI5/MM842_g N_VSS_XI5/MM842_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1479 XI5/NET01770 N_NET38_XI5/MM1479_g N_VSS_XI5/MM1479_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM821 N_NET160_XI5/MM821_d N_NET39_XI5/MM821_g N_VSS_XI5/MM821_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1471 XI5/NET01802 N_NET40_XI5/MM1471_g N_VSS_XI5/MM1471_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM810 N_NET160_XI5/MM810_d N_NET41_XI5/MM810_g N_VSS_XI5/MM810_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1463 XI5/NET01834 N_NET42_XI5/MM1463_g N_VSS_XI5/MM1463_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM789 N_NET160_XI5/MM789_d N_NET43_XI5/MM789_g N_VSS_XI5/MM789_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1455 XI5/NET01866 N_NET44_XI5/MM1455_g N_VSS_XI5/MM1455_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM778 N_NET160_XI5/MM778_d N_NET45_XI5/MM778_g N_VSS_XI5/MM778_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1447 XI5/NET01898 N_NET46_XI5/MM1447_g N_VSS_XI5/MM1447_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM757 N_NET160_XI5/MM757_d N_NET47_XI5/MM757_g N_VSS_XI5/MM757_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1439 XI5/NET01930 N_NET48_XI5/MM1439_g N_VSS_XI5/MM1439_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM746 N_NET160_XI5/MM746_d N_NET49_XI5/MM746_g N_VSS_XI5/MM746_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1431 XI5/NET01962 N_NET50_XI5/MM1431_g N_VSS_XI5/MM1431_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM730 N_NET160_XI5/MM730_d N_NET51_XI5/MM730_g N_VSS_XI5/MM730_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1423 XI5/NET01994 N_NET52_XI5/MM1423_g N_VSS_XI5/MM1423_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM709 N_NET160_XI5/MM709_d N_NET53_XI5/MM709_g N_VSS_XI5/MM709_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1415 XI5/NET02026 N_NET54_XI5/MM1415_g N_VSS_XI5/MM1415_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM698 N_NET160_XI5/MM698_d N_NET55_XI5/MM698_g N_VSS_XI5/MM698_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1407 XI5/NET02058 N_NET56_XI5/MM1407_g N_VSS_XI5/MM1407_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM677 N_NET160_XI5/MM677_d N_NET57_XI5/MM677_g N_VSS_XI5/MM677_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1399 XI5/NET02090 N_NET58_XI5/MM1399_g N_VSS_XI5/MM1399_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM666 N_NET160_XI5/MM666_d N_NET59_XI5/MM666_g N_VSS_XI5/MM666_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1391 XI5/NET02122 N_NET60_XI5/MM1391_g N_VSS_XI5/MM1391_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM645 N_NET160_XI5/MM645_d N_NET61_XI5/MM645_g N_VSS_XI5/MM645_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1383 XI5/NET02154 N_NET62_XI5/MM1383_g N_VSS_XI5/MM1383_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM634 N_NET160_XI5/MM634_d N_NET63_XI5/MM634_g N_VSS_XI5/MM634_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1375 XI5/NET02186 N_NET64_XI5/MM1375_g N_VSS_XI5/MM1375_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM613 N_NET160_XI5/MM613_d N_NET65_XI5/MM613_g N_VSS_XI5/MM613_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1367 XI5/NET02218 N_NET66_XI5/MM1367_g N_VSS_XI5/MM1367_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM596 N_NET160_XI5/MM596_d N_NET67_XI5/MM596_g N_VSS_XI5/MM596_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1359 XI5/NET02250 N_NET68_XI5/MM1359_g N_VSS_XI5/MM1359_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM587 N_NET160_XI5/MM587_d N_NET69_XI5/MM587_g N_VSS_XI5/MM587_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1347 XI5/NET02298 N_NET70_XI5/MM1347_g N_VSS_XI5/MM1347_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM541 N_NET160_XI5/MM541_d N_NET71_XI5/MM541_g N_VSS_XI5/MM541_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1065 XI5/NET04434 N_NET72_XI5/MM1065_g N_VSS_XI5/MM1065_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM521 N_NET160_XI5/MM521_d N_NET8_XI5/MM521_g N_VSS_XI5/MM521_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM37 N_XI7/NET45_XI7/MM37_d N_NET125_XI7/MM37_g N_XI7/NET69_XI7/MM37_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI7/MM36 N_XI7/NET49_XI7/MM36_d N_XI7/NET68_XI7/MM36_g N_XI7/NET69_XI7/MM36_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI7/MM40 N_NET161_XI7/MM40_d N_NET120_XI7/MM40_g N_XI7/NET49_XI7/MM40_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI5/MM1049 N_NET161_XI5/MM1049_d N_NET10_XI5/MM1049_g N_VSS_XI5/MM1049_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1330 XI5/NET02334 N_NET11_XI5/MM1330_g N_VSS_XI5/MM1330_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1030 N_NET161_XI5/MM1030_d N_NET12_XI5/MM1030_g N_VSS_XI5/MM1030_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1328 XI5/NET02342 N_NET13_XI5/MM1328_g N_VSS_XI5/MM1328_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1017 N_NET161_XI5/MM1017_d N_NET14_XI5/MM1017_g N_VSS_XI5/MM1017_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1320 XI5/NET02374 N_NET15_XI5/MM1320_g N_VSS_XI5/MM1320_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM998 N_NET161_XI5/MM998_d N_NET16_XI5/MM998_g N_VSS_XI5/MM998_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1312 XI5/NET02406 N_NET17_XI5/MM1312_g N_VSS_XI5/MM1312_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM985 N_NET161_XI5/MM985_d N_NET18_XI5/MM985_g N_VSS_XI5/MM985_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1304 XI5/NET02438 N_NET19_XI5/MM1304_g N_VSS_XI5/MM1304_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM966 N_NET161_XI5/MM966_d N_NET20_XI5/MM966_g N_VSS_XI5/MM966_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1296 XI5/NET04258 N_NET21_XI5/MM1296_g N_VSS_XI5/MM1296_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM953 N_NET161_XI5/MM953_d N_NET22_XI5/MM953_g N_VSS_XI5/MM953_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1288 XI5/NET04290 N_NET23_XI5/MM1288_g N_VSS_XI5/MM1288_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM934 N_NET161_XI5/MM934_d N_NET24_XI5/MM934_g N_VSS_XI5/MM934_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1280 XI5/NET03438 N_NET25_XI5/MM1280_g N_VSS_XI5/MM1280_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM921 N_NET161_XI5/MM921_d N_NET26_XI5/MM921_g N_VSS_XI5/MM921_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1265 XI5/NET05378 N_NET27_XI5/MM1265_g N_VSS_XI5/MM1265_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM902 N_NET161_XI5/MM902_d N_NET28_XI5/MM902_g N_VSS_XI5/MM902_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1257 XI5/NET05334 N_NET29_XI5/MM1257_g N_VSS_XI5/MM1257_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM889 N_NET161_XI5/MM889_d N_NET30_XI5/MM889_g N_VSS_XI5/MM889_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1249 XI5/NET05290 N_NET31_XI5/MM1249_g N_VSS_XI5/MM1249_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM870 N_NET161_XI5/MM870_d N_NET32_XI5/MM870_g N_VSS_XI5/MM870_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1241 XI5/NET05258 N_NET33_XI5/MM1241_g N_VSS_XI5/MM1241_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM857 N_NET161_XI5/MM857_d N_NET34_XI5/MM857_g N_VSS_XI5/MM857_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1233 XI5/NET05226 N_NET35_XI5/MM1233_g N_VSS_XI5/MM1233_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM838 N_NET161_XI5/MM838_d N_NET36_XI5/MM838_g N_VSS_XI5/MM838_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1225 XI5/NET05194 N_NET37_XI5/MM1225_g N_VSS_XI5/MM1225_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM825 N_NET161_XI5/MM825_d N_NET38_XI5/MM825_g N_VSS_XI5/MM825_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1217 XI5/NET05154 N_NET39_XI5/MM1217_g N_VSS_XI5/MM1217_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM806 N_NET161_XI5/MM806_d N_NET40_XI5/MM806_g N_VSS_XI5/MM806_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1209 XI5/NET05122 N_NET41_XI5/MM1209_g N_VSS_XI5/MM1209_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM793 N_NET161_XI5/MM793_d N_NET42_XI5/MM793_g N_VSS_XI5/MM793_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1201 XI5/NET05086 N_NET43_XI5/MM1201_g N_VSS_XI5/MM1201_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM774 N_NET161_XI5/MM774_d N_NET44_XI5/MM774_g N_VSS_XI5/MM774_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1193 XI5/NET05054 N_NET45_XI5/MM1193_g N_VSS_XI5/MM1193_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM761 N_NET161_XI5/MM761_d N_NET46_XI5/MM761_g N_VSS_XI5/MM761_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1185 XI5/NET05022 N_NET47_XI5/MM1185_g N_VSS_XI5/MM1185_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM742 N_NET161_XI5/MM742_d N_NET48_XI5/MM742_g N_VSS_XI5/MM742_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1177 XI5/NET04990 N_NET49_XI5/MM1177_g N_VSS_XI5/MM1177_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM726 N_NET161_XI5/MM726_d N_NET50_XI5/MM726_g N_VSS_XI5/MM726_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1169 XI5/NET04958 N_NET51_XI5/MM1169_g N_VSS_XI5/MM1169_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM713 N_NET161_XI5/MM713_d N_NET52_XI5/MM713_g N_VSS_XI5/MM713_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1161 XI5/NET04926 N_NET53_XI5/MM1161_g N_VSS_XI5/MM1161_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM694 N_NET161_XI5/MM694_d N_NET54_XI5/MM694_g N_VSS_XI5/MM694_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1153 XI5/NET04886 N_NET55_XI5/MM1153_g N_VSS_XI5/MM1153_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM681 N_NET161_XI5/MM681_d N_NET56_XI5/MM681_g N_VSS_XI5/MM681_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1145 XI5/NET04854 N_NET57_XI5/MM1145_g N_VSS_XI5/MM1145_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM662 N_NET161_XI5/MM662_d N_NET58_XI5/MM662_g N_VSS_XI5/MM662_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1137 XI5/NET04822 N_NET59_XI5/MM1137_g N_VSS_XI5/MM1137_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM649 N_NET161_XI5/MM649_d N_NET60_XI5/MM649_g N_VSS_XI5/MM649_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1129 XI5/NET04790 N_NET61_XI5/MM1129_g N_VSS_XI5/MM1129_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM630 N_NET161_XI5/MM630_d N_NET62_XI5/MM630_g N_VSS_XI5/MM630_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1122 XI5/NET04738 N_NET63_XI5/MM1122_g N_VSS_XI5/MM1122_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM617 N_NET161_XI5/MM617_d N_NET64_XI5/MM617_g N_VSS_XI5/MM617_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1097 XI5/NET04666 N_NET65_XI5/MM1097_g N_VSS_XI5/MM1097_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM600 N_NET161_XI5/MM600_d N_NET66_XI5/MM600_g N_VSS_XI5/MM600_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1088 XI5/NET04622 N_NET67_XI5/MM1088_g N_VSS_XI5/MM1088_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM583 N_NET161_XI5/MM583_d N_NET68_XI5/MM583_g N_VSS_XI5/MM583_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1080 XI5/NET04590 N_NET69_XI5/MM1080_g N_VSS_XI5/MM1080_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM531 N_NET161_XI5/MM531_d N_NET70_XI5/MM531_g N_VSS_XI5/MM531_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1072 XI5/NET04546 N_NET71_XI5/MM1072_g N_VSS_XI5/MM1072_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM528 N_NET161_XI5/MM528_d N_NET72_XI5/MM528_g N_VSS_XI5/MM528_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1056 XI5/NET02746 N_NET8_XI5/MM1056_g N_VSS_XI5/MM1056_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM41 N_NET162_XI7/MM41_d N_XI7/NET48_XI7/MM41_g N_XI7/NET49_XI7/MM41_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXI5/MM1592 XI5/NET01318 N_NET10_XI5/MM1592_g N_VSS_XI5/MM1592_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1042 N_NET162_XI5/MM1042_d N_NET11_XI5/MM1042_g N_VSS_XI5/MM1042_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1584 XI5/NET01350 N_NET12_XI5/MM1584_g N_VSS_XI5/MM1584_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1037 N_NET162_XI5/MM1037_d N_NET13_XI5/MM1037_g N_VSS_XI5/MM1037_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1576 XI5/NET01382 N_NET14_XI5/MM1576_g N_VSS_XI5/MM1576_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1010 N_NET162_XI5/MM1010_d N_NET15_XI5/MM1010_g N_VSS_XI5/MM1010_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1568 XI5/NET01414 N_NET16_XI5/MM1568_g N_VSS_XI5/MM1568_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1005 N_NET162_XI5/MM1005_d N_NET17_XI5/MM1005_g N_VSS_XI5/MM1005_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1560 XI5/NET01446 N_NET18_XI5/MM1560_g N_VSS_XI5/MM1560_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM978 N_NET162_XI5/MM978_d N_NET19_XI5/MM978_g N_VSS_XI5/MM978_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1552 XI5/NET01478 N_NET20_XI5/MM1552_g N_VSS_XI5/MM1552_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM973 N_NET162_XI5/MM973_d N_NET21_XI5/MM973_g N_VSS_XI5/MM973_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1544 XI5/NET01510 N_NET22_XI5/MM1544_g N_VSS_XI5/MM1544_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM946 N_NET162_XI5/MM946_d N_NET23_XI5/MM946_g N_VSS_XI5/MM946_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1536 XI5/NET01542 N_NET24_XI5/MM1536_g N_VSS_XI5/MM1536_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM941 N_NET162_XI5/MM941_d N_NET25_XI5/MM941_g N_VSS_XI5/MM941_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1528 XI5/NET01574 N_NET26_XI5/MM1528_g N_VSS_XI5/MM1528_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM914 N_NET162_XI5/MM914_d N_NET27_XI5/MM914_g N_VSS_XI5/MM914_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1520 XI5/NET01606 N_NET28_XI5/MM1520_g N_VSS_XI5/MM1520_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM909 N_NET162_XI5/MM909_d N_NET29_XI5/MM909_g N_VSS_XI5/MM909_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1512 XI5/NET01638 N_NET30_XI5/MM1512_g N_VSS_XI5/MM1512_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM882 N_NET162_XI5/MM882_d N_NET31_XI5/MM882_g N_VSS_XI5/MM882_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1504 XI5/NET01670 N_NET32_XI5/MM1504_g N_VSS_XI5/MM1504_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM877 N_NET162_XI5/MM877_d N_NET33_XI5/MM877_g N_VSS_XI5/MM877_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1496 XI5/NET01702 N_NET34_XI5/MM1496_g N_VSS_XI5/MM1496_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM850 N_NET162_XI5/MM850_d N_NET35_XI5/MM850_g N_VSS_XI5/MM850_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1488 XI5/NET01734 N_NET36_XI5/MM1488_g N_VSS_XI5/MM1488_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM845 N_NET162_XI5/MM845_d N_NET37_XI5/MM845_g N_VSS_XI5/MM845_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1480 XI5/NET01766 N_NET38_XI5/MM1480_g N_VSS_XI5/MM1480_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM818 N_NET162_XI5/MM818_d N_NET39_XI5/MM818_g N_VSS_XI5/MM818_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1472 XI5/NET01798 N_NET40_XI5/MM1472_g N_VSS_XI5/MM1472_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM813 N_NET162_XI5/MM813_d N_NET41_XI5/MM813_g N_VSS_XI5/MM813_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1464 XI5/NET01830 N_NET42_XI5/MM1464_g N_VSS_XI5/MM1464_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM786 N_NET162_XI5/MM786_d N_NET43_XI5/MM786_g N_VSS_XI5/MM786_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1456 XI5/NET01862 N_NET44_XI5/MM1456_g N_VSS_XI5/MM1456_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM781 N_NET162_XI5/MM781_d N_NET45_XI5/MM781_g N_VSS_XI5/MM781_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1448 XI5/NET01894 N_NET46_XI5/MM1448_g N_VSS_XI5/MM1448_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM754 N_NET162_XI5/MM754_d N_NET47_XI5/MM754_g N_VSS_XI5/MM754_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1440 XI5/NET01926 N_NET48_XI5/MM1440_g N_VSS_XI5/MM1440_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM749 N_NET162_XI5/MM749_d N_NET49_XI5/MM749_g N_VSS_XI5/MM749_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1432 XI5/NET01958 N_NET50_XI5/MM1432_g N_VSS_XI5/MM1432_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM733 N_NET162_XI5/MM733_d N_NET51_XI5/MM733_g N_VSS_XI5/MM733_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1424 XI5/NET01990 N_NET52_XI5/MM1424_g N_VSS_XI5/MM1424_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM706 N_NET162_XI5/MM706_d N_NET53_XI5/MM706_g N_VSS_XI5/MM706_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1416 XI5/NET02022 N_NET54_XI5/MM1416_g N_VSS_XI5/MM1416_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM701 N_NET162_XI5/MM701_d N_NET55_XI5/MM701_g N_VSS_XI5/MM701_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1408 XI5/NET02054 N_NET56_XI5/MM1408_g N_VSS_XI5/MM1408_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM674 N_NET162_XI5/MM674_d N_NET57_XI5/MM674_g N_VSS_XI5/MM674_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1400 XI5/NET02086 N_NET58_XI5/MM1400_g N_VSS_XI5/MM1400_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM669 N_NET162_XI5/MM669_d N_NET59_XI5/MM669_g N_VSS_XI5/MM669_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1392 XI5/NET02118 N_NET60_XI5/MM1392_g N_VSS_XI5/MM1392_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM642 N_NET162_XI5/MM642_d N_NET61_XI5/MM642_g N_VSS_XI5/MM642_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1384 XI5/NET02150 N_NET62_XI5/MM1384_g N_VSS_XI5/MM1384_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM637 N_NET162_XI5/MM637_d N_NET63_XI5/MM637_g N_VSS_XI5/MM637_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1376 XI5/NET02182 N_NET64_XI5/MM1376_g N_VSS_XI5/MM1376_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM610 N_NET162_XI5/MM610_d N_NET65_XI5/MM610_g N_VSS_XI5/MM610_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1368 XI5/NET02214 N_NET66_XI5/MM1368_g N_VSS_XI5/MM1368_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM593 N_NET162_XI5/MM593_d N_NET67_XI5/MM593_g N_VSS_XI5/MM593_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1360 XI5/NET02246 N_NET68_XI5/MM1360_g N_VSS_XI5/MM1360_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM590 N_NET162_XI5/MM590_d N_NET69_XI5/MM590_g N_VSS_XI5/MM590_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1346 XI5/NET02302 N_NET70_XI5/MM1346_g N_VSS_XI5/MM1346_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM544 N_NET162_XI5/MM544_d N_NET71_XI5/MM544_g N_VSS_XI5/MM544_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM1064 XI5/NET04394 N_NET72_XI5/MM1064_g N_VSS_XI5/MM1064_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI5/MM520 N_NET162_XI5/MM520_d N_NET8_XI5/MM520_g N_VSS_XI5/MM520_s
+ N_VSS_XI45/XI0/XI8/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI45/XI0/XI8/MM1 N_XI45/XI0/NET96_XI45/XI0/XI8/MM1_d
+ N_NET100_XI45/XI0/XI8/MM1_g N_VDD_XI45/XI0/XI8/MM1_s N_VDD_XI45/XI0/XI8/MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI45/XI1/XI8/MM1 N_XI45/XI1/NET96_XI45/XI1/XI8/MM1_d
+ N_NET110_XI45/XI1/XI8/MM1_g N_VDD_XI45/XI1/XI8/MM1_s N_VDD_XI45/XI0/XI8/MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI45/XI0/XI9/MM1 N_XI45/XI0/NET92_XI45/XI0/XI9/MM1_d
+ N_NET105_XI45/XI0/XI9/MM1_g N_VDD_XI45/XI0/XI9/MM1_s N_VDD_XI45/XI0/XI8/MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI45/XI1/XI9/MM1 N_XI45/XI1/NET92_XI45/XI1/XI9/MM1_d N_NET90_XI45/XI1/XI9/MM1_g
+ N_VDD_XI45/XI1/XI9/MM1_s N_VDD_XI45/XI0/XI8/MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI46/MM4 N_DOUT<1>_XI46/MM4_d N_NET0176_XI46/MM4_g N_VDD_XI46/MM4_s
+ N_VDD_XI46/MM4_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=3.6e-13 PD=1.98e-06
+ PS=7.2e-07
mXI46/MM5 N_NET0176_XI46/MM5_d N_DOUT<1>_XI46/MM5_g N_VDD_XI46/MM5_s
+ N_VDD_XI46/MM4_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=3.6e-13 PD=1.98e-06
+ PS=7.2e-07
mXI10/MM0 N_XI10/NET28_XI10/MM0_d N_A<7>_XI10/MM0_g N_VDD_XI10/MM0_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=1.875e-13 AS=7.35e-13 PD=2.5e-07
+ PS=2.48e-06
mXI10/MM4 N_XI10/NET13_XI10/MM4_d N_CLK_XI10/MM4_g N_XI10/NET28_XI10/MM4_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=1.875e-13 PD=2.48e-06
+ PS=2.5e-07
mXI10/MM1 N_XI10/NET21_XI10/MM1_d N_CLK_XI10/MM1_g N_VDD_XI10/MM1_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI10/MM2 N_XI10/NET15_XI10/MM2_d N_XI10/NET21_XI10/MM2_g N_VDD_XI10/MM2_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=6.11842e-13 AS=7.35e-13
+ PD=1.8e-06 PS=2.48e-06
mXI10/MM3 N_NET125_XI10/MM3_d N_XI10/NET15_XI10/MM3_g N_VDD_XI10/MM3_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=6.11842e-13
+ PD=2.48e-06 PS=1.8e-06
mXI18/MM0 N_XI18/NET28_XI18/MM0_d N_A<6>_XI18/MM0_g N_VDD_XI18/MM0_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=1.875e-13 AS=7.35e-13 PD=2.5e-07
+ PS=2.48e-06
mXI18/MM4 N_XI18/NET13_XI18/MM4_d N_CLK_XI18/MM4_g N_XI18/NET28_XI18/MM4_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=1.875e-13 PD=2.48e-06
+ PS=2.5e-07
mXI18/MM1 N_XI18/NET21_XI18/MM1_d N_CLK_XI18/MM1_g N_VDD_XI18/MM1_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI18/MM2 N_XI18/NET15_XI18/MM2_d N_XI18/NET21_XI18/MM2_g N_VDD_XI18/MM2_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=6.11842e-13 AS=7.35e-13
+ PD=1.8e-06 PS=2.48e-06
mXI18/MM3 N_NET85_XI18/MM3_d N_XI18/NET15_XI18/MM3_g N_VDD_XI18/MM3_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=6.11842e-13
+ PD=2.48e-06 PS=1.8e-06
mXI16/MM0 N_XI16/NET28_XI16/MM0_d N_A<2>_XI16/MM0_g N_VDD_XI16/MM0_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=1.875e-13 AS=7.35e-13 PD=2.5e-07
+ PS=2.48e-06
mXI16/MM4 N_XI16/NET13_XI16/MM4_d N_CLK_XI16/MM4_g N_XI16/NET28_XI16/MM4_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=1.875e-13 PD=2.48e-06
+ PS=2.5e-07
mXI16/MM1 N_XI16/NET21_XI16/MM1_d N_CLK_XI16/MM1_g N_VDD_XI16/MM1_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI16/MM2 N_XI16/NET15_XI16/MM2_d N_XI16/NET21_XI16/MM2_g N_VDD_XI16/MM2_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=6.11842e-13 AS=7.35e-13
+ PD=1.8e-06 PS=2.48e-06
mXI16/MM3 N_NET95_XI16/MM3_d N_XI16/NET15_XI16/MM3_g N_VDD_XI16/MM3_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=6.11842e-13
+ PD=2.48e-06 PS=1.8e-06
mXI14/MM0 N_XI14/NET28_XI14/MM0_d N_A<1>_XI14/MM0_g N_VDD_XI14/MM0_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=1.875e-13 AS=7.35e-13 PD=2.5e-07
+ PS=2.48e-06
mXI14/MM4 N_XI14/NET13_XI14/MM4_d N_CLK_XI14/MM4_g N_XI14/NET28_XI14/MM4_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=1.875e-13 PD=2.48e-06
+ PS=2.5e-07
mXI14/MM1 N_XI14/NET21_XI14/MM1_d N_CLK_XI14/MM1_g N_VDD_XI14/MM1_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI14/MM2 N_XI14/NET15_XI14/MM2_d N_XI14/NET21_XI14/MM2_g N_VDD_XI14/MM2_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=6.11842e-13 AS=7.35e-13
+ PD=1.8e-06 PS=2.48e-06
mXI14/MM3 N_NET105_XI14/MM3_d N_XI14/NET15_XI14/MM3_g N_VDD_XI14/MM3_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=6.11842e-13
+ PD=2.48e-06 PS=1.8e-06
mXI15/MM0 N_XI15/NET28_XI15/MM0_d N_A<0>_XI15/MM0_g N_VDD_XI15/MM0_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=1.875e-13 AS=7.35e-13 PD=2.5e-07
+ PS=2.48e-06
mXI15/MM4 N_XI15/NET13_XI15/MM4_d N_CLK_XI15/MM4_g N_XI15/NET28_XI15/MM4_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=1.875e-13 PD=2.48e-06
+ PS=2.5e-07
mXI15/MM1 N_XI15/NET21_XI15/MM1_d N_CLK_XI15/MM1_g N_VDD_XI15/MM1_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15/MM2 N_XI15/NET15_XI15/MM2_d N_XI15/NET21_XI15/MM2_g N_VDD_XI15/MM2_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=6.11842e-13 AS=7.35e-13
+ PD=1.8e-06 PS=2.48e-06
mXI15/MM3 N_NET100_XI15/MM3_d N_XI15/NET15_XI15/MM3_g N_VDD_XI15/MM3_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=6.11842e-13
+ PD=2.48e-06 PS=1.8e-06
mXI45/XI0/XI10/MM1 N_XI45/XI0/NET081_XI45/XI0/XI10/MM1_d
+ N_NET95_XI45/XI0/XI10/MM1_g N_VDD_XI45/XI0/XI10/MM1_s N_VDD_XI45/XI0/XI8/MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI45/XI1/XI10/MM1 N_XI45/XI1/NET081_XI45/XI1/XI10/MM1_d
+ N_NET115_XI45/XI1/XI10/MM1_g N_VDD_XI45/XI1/XI10/MM1_s
+ N_VDD_XI45/XI0/XI8/MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI10/MM11 N_XI10/NET15_XI10/MM11_d N_NET125_XI10/MM11_g N_VDD_XI10/MM11_s
+ N_VDD_XI10/MM0_b P_18 L=5.3e-07 W=4e-07 AD=1.63158e-13 AS=1.63158e-13
+ PD=4.8e-07 PS=4.8e-07
mXI18/MM11 N_XI18/NET15_XI18/MM11_d N_NET85_XI18/MM11_g N_VDD_XI18/MM11_s
+ N_VDD_XI10/MM0_b P_18 L=5.3e-07 W=4e-07 AD=1.63158e-13 AS=1.63158e-13
+ PD=4.8e-07 PS=4.8e-07
mXI16/MM11 N_XI16/NET15_XI16/MM11_d N_NET95_XI16/MM11_g N_VDD_XI16/MM11_s
+ N_VDD_XI10/MM0_b P_18 L=5.3e-07 W=4e-07 AD=1.63158e-13 AS=1.63158e-13
+ PD=4.8e-07 PS=4.8e-07
mXI14/MM11 N_XI14/NET15_XI14/MM11_d N_NET105_XI14/MM11_g N_VDD_XI14/MM11_s
+ N_VDD_XI10/MM0_b P_18 L=5.3e-07 W=4e-07 AD=1.63158e-13 AS=1.63158e-13
+ PD=4.8e-07 PS=4.8e-07
mXI15/MM11 N_XI15/NET15_XI15/MM11_d N_NET100_XI15/MM11_g N_VDD_XI15/MM11_s
+ N_VDD_XI10/MM0_b P_18 L=5.3e-07 W=4e-07 AD=1.63158e-13 AS=1.63158e-13
+ PD=4.8e-07 PS=4.8e-07
mXI19/MM6 N_XI19/NET0139_XI19/MM6_d N_XI19/NET41_XI19/MM6_g N_VDD_XI19/MM6_s
+ N_VDD_XI10/MM0_b P_18 L=8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI19/MM5 N_XI19/NET41_XI19/MM5_d N_CLK_XI19/MM5_g N_VDD_XI19/MM5_s
+ N_VDD_XI10/MM0_b P_18 L=8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI19/MM3 N_NET81_XI19/MM3_d N_XI19/NET49_XI19/MM3_g N_VDD_XI19/MM3_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI19/MM0 N_XI19/NET49_XI19/MM0_d N_CLK_XI19/MM0_g N_VDD_XI19/MM0_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI11/MM0 N_XI11/NET28_XI11/MM0_d N_A<8>_XI11/MM0_g N_VDD_XI11/MM0_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=1.875e-13 AS=7.35e-13 PD=2.5e-07
+ PS=2.48e-06
mXI11/MM4 N_XI11/NET13_XI11/MM4_d N_CLK_XI11/MM4_g N_XI11/NET28_XI11/MM4_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=1.875e-13 PD=2.48e-06
+ PS=2.5e-07
mXI11/MM1 N_XI11/NET21_XI11/MM1_d N_CLK_XI11/MM1_g N_VDD_XI11/MM1_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI11/MM2 N_XI11/NET15_XI11/MM2_d N_XI11/NET21_XI11/MM2_g N_VDD_XI11/MM2_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=6.11842e-13 AS=7.35e-13
+ PD=1.8e-06 PS=2.48e-06
mXI11/MM11 N_XI11/NET15_XI11/MM11_d N_NET120_XI11/MM11_g N_VDD_XI11/MM11_s
+ N_VDD_XI10/MM0_b P_18 L=5.3e-07 W=4e-07 AD=1.63158e-13 AS=1.63158e-13
+ PD=4.8e-07 PS=4.8e-07
mXI11/MM3 N_NET120_XI11/MM3_d N_XI11/NET15_XI11/MM3_g N_VDD_XI11/MM3_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=6.11842e-13
+ PD=2.48e-06 PS=1.8e-06
mXI12/MM0 N_XI12/NET28_XI12/MM0_d N_A<5>_XI12/MM0_g N_VDD_XI12/MM0_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=1.875e-13 AS=7.35e-13 PD=2.5e-07
+ PS=2.48e-06
mXI12/MM4 N_XI12/NET13_XI12/MM4_d N_CLK_XI12/MM4_g N_XI12/NET28_XI12/MM4_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=1.875e-13 PD=2.48e-06
+ PS=2.5e-07
mXI12/MM1 N_XI12/NET21_XI12/MM1_d N_CLK_XI12/MM1_g N_VDD_XI12/MM1_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI12/MM2 N_XI12/NET15_XI12/MM2_d N_XI12/NET21_XI12/MM2_g N_VDD_XI12/MM2_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=6.11842e-13 AS=7.35e-13
+ PD=1.8e-06 PS=2.48e-06
mXI12/MM11 N_XI12/NET15_XI12/MM11_d N_NET115_XI12/MM11_g N_VDD_XI12/MM11_s
+ N_VDD_XI10/MM0_b P_18 L=5.3e-07 W=4e-07 AD=1.63158e-13 AS=1.63158e-13
+ PD=4.8e-07 PS=4.8e-07
mXI12/MM3 N_NET115_XI12/MM3_d N_XI12/NET15_XI12/MM3_g N_VDD_XI12/MM3_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=6.11842e-13
+ PD=2.48e-06 PS=1.8e-06
mXI17/MM0 N_XI17/NET28_XI17/MM0_d N_A<4>_XI17/MM0_g N_VDD_XI17/MM0_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=1.875e-13 AS=7.35e-13 PD=2.5e-07
+ PS=2.48e-06
mXI17/MM4 N_XI17/NET13_XI17/MM4_d N_CLK_XI17/MM4_g N_XI17/NET28_XI17/MM4_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=1.875e-13 PD=2.48e-06
+ PS=2.5e-07
mXI17/MM1 N_XI17/NET21_XI17/MM1_d N_CLK_XI17/MM1_g N_VDD_XI17/MM1_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI17/MM2 N_XI17/NET15_XI17/MM2_d N_XI17/NET21_XI17/MM2_g N_VDD_XI17/MM2_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=6.11842e-13 AS=7.35e-13
+ PD=1.8e-06 PS=2.48e-06
mXI17/MM11 N_XI17/NET15_XI17/MM11_d N_NET90_XI17/MM11_g N_VDD_XI17/MM11_s
+ N_VDD_XI10/MM0_b P_18 L=5.3e-07 W=4e-07 AD=1.63158e-13 AS=1.63158e-13
+ PD=4.8e-07 PS=4.8e-07
mXI17/MM3 N_NET90_XI17/MM3_d N_XI17/NET15_XI17/MM3_g N_VDD_XI17/MM3_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=6.11842e-13
+ PD=2.48e-06 PS=1.8e-06
mXI13/MM0 N_XI13/NET28_XI13/MM0_d N_A<3>_XI13/MM0_g N_VDD_XI13/MM0_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=1.875e-13 AS=7.35e-13 PD=2.5e-07
+ PS=2.48e-06
mXI13/MM4 N_XI13/NET13_XI13/MM4_d N_CLK_XI13/MM4_g N_XI13/NET28_XI13/MM4_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=1.875e-13 PD=2.48e-06
+ PS=2.5e-07
mXI13/MM1 N_XI13/NET21_XI13/MM1_d N_CLK_XI13/MM1_g N_VDD_XI13/MM1_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI13/MM2 N_XI13/NET15_XI13/MM2_d N_XI13/NET21_XI13/MM2_g N_VDD_XI13/MM2_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=6.11842e-13 AS=7.35e-13
+ PD=1.8e-06 PS=2.48e-06
mXI13/MM11 N_XI13/NET15_XI13/MM11_d N_NET110_XI13/MM11_g N_VDD_XI13/MM11_s
+ N_VDD_XI10/MM0_b P_18 L=5.3e-07 W=4e-07 AD=1.63158e-13 AS=1.63158e-13
+ PD=4.8e-07 PS=4.8e-07
mXI13/MM3 N_NET110_XI13/MM3_d N_XI13/NET15_XI13/MM3_g N_VDD_XI13/MM3_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=6.11842e-13
+ PD=2.48e-06 PS=1.8e-06
mXI47/MM4 N_DOUT<0>_XI47/MM4_d N_NET0183_XI47/MM4_g N_VDD_XI47/MM4_s
+ N_VDD_XI46/MM4_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=3.6e-13 PD=1.98e-06
+ PS=7.2e-07
mXI47/MM5 N_NET0183_XI47/MM5_d N_DOUT<0>_XI47/MM5_g N_VDD_XI47/MM5_s
+ N_VDD_XI46/MM4_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=3.6e-13 PD=1.98e-06
+ PS=7.2e-07
mXI45/XI0/XI18/MM3 N_XI45/NET272_XI45/XI0/XI18/MM3_d N_NET79_XI45/XI0/XI18/MM3_g
+ N_VDD_XI45/XI0/XI18/MM3_s N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI18/MM2 N_XI45/NET272_XI45/XI0/XI18/MM2_d
+ N_XI45/XI0/NET081_XI45/XI0/XI18/MM2_g N_VDD_XI45/XI0/XI18/MM2_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07
+ PS=5.4e-07
mXI45/XI0/XI18/MM1 N_XI45/NET272_XI45/XI0/XI18/MM1_d
+ N_XI45/XI0/NET92_XI45/XI0/XI18/MM1_g N_VDD_XI45/XI0/XI18/MM1_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07
+ PS=5.4e-07
mXI45/XI0/XI18/MM0 N_XI45/NET272_XI45/XI0/XI18/MM0_d
+ N_XI45/XI0/NET96_XI45/XI0/XI18/MM0_g N_VDD_XI45/XI0/XI18/MM0_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13
+ PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI17/MM3 N_XI45/NET273_XI45/XI0/XI17/MM3_d N_NET79_XI45/XI0/XI17/MM3_g
+ N_VDD_XI45/XI0/XI17/MM3_s N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI17/MM2 N_XI45/NET273_XI45/XI0/XI17/MM2_d N_NET95_XI45/XI0/XI17/MM2_g
+ N_VDD_XI45/XI0/XI17/MM2_s N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI17/MM1 N_XI45/NET273_XI45/XI0/XI17/MM1_d
+ N_XI45/XI0/NET92_XI45/XI0/XI17/MM1_g N_VDD_XI45/XI0/XI17/MM1_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07
+ PS=5.4e-07
mXI45/XI0/XI17/MM0 N_XI45/NET273_XI45/XI0/XI17/MM0_d
+ N_XI45/XI0/NET96_XI45/XI0/XI17/MM0_g N_VDD_XI45/XI0/XI17/MM0_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13
+ PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI16/MM3 N_XI45/NET274_XI45/XI0/XI16/MM3_d N_NET79_XI45/XI0/XI16/MM3_g
+ N_VDD_XI45/XI0/XI16/MM3_s N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI16/MM2 N_XI45/NET274_XI45/XI0/XI16/MM2_d
+ N_XI45/XI0/NET081_XI45/XI0/XI16/MM2_g N_VDD_XI45/XI0/XI16/MM2_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07
+ PS=5.4e-07
mXI45/XI0/XI16/MM1 N_XI45/NET274_XI45/XI0/XI16/MM1_d
+ N_NET105_XI45/XI0/XI16/MM1_g N_VDD_XI45/XI0/XI16/MM1_s N_VDD_XI10/MM0_b P_18
+ L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI16/MM0 N_XI45/NET274_XI45/XI0/XI16/MM0_d
+ N_XI45/XI0/NET96_XI45/XI0/XI16/MM0_g N_VDD_XI45/XI0/XI16/MM0_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13
+ PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI15/MM3 N_XI45/NET275_XI45/XI0/XI15/MM3_d N_NET79_XI45/XI0/XI15/MM3_g
+ N_VDD_XI45/XI0/XI15/MM3_s N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI15/MM2 N_XI45/NET275_XI45/XI0/XI15/MM2_d N_NET95_XI45/XI0/XI15/MM2_g
+ N_VDD_XI45/XI0/XI15/MM2_s N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI15/MM1 N_XI45/NET275_XI45/XI0/XI15/MM1_d
+ N_NET105_XI45/XI0/XI15/MM1_g N_VDD_XI45/XI0/XI15/MM1_s N_VDD_XI10/MM0_b P_18
+ L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI15/MM0 N_XI45/NET275_XI45/XI0/XI15/MM0_d
+ N_XI45/XI0/NET96_XI45/XI0/XI15/MM0_g N_VDD_XI45/XI0/XI15/MM0_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13
+ PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI14/MM3 N_XI45/NET276_XI45/XI0/XI14/MM3_d N_NET79_XI45/XI0/XI14/MM3_g
+ N_VDD_XI45/XI0/XI14/MM3_s N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI14/MM2 N_XI45/NET276_XI45/XI0/XI14/MM2_d
+ N_XI45/XI0/NET081_XI45/XI0/XI14/MM2_g N_VDD_XI45/XI0/XI14/MM2_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07
+ PS=5.4e-07
mXI45/XI0/XI14/MM1 N_XI45/NET276_XI45/XI0/XI14/MM1_d
+ N_XI45/XI0/NET92_XI45/XI0/XI14/MM1_g N_VDD_XI45/XI0/XI14/MM1_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07
+ PS=5.4e-07
mXI45/XI0/XI14/MM0 N_XI45/NET276_XI45/XI0/XI14/MM0_d
+ N_NET100_XI45/XI0/XI14/MM0_g N_VDD_XI45/XI0/XI14/MM0_s N_VDD_XI10/MM0_b P_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI13/MM3 N_XI45/NET277_XI45/XI0/XI13/MM3_d N_NET79_XI45/XI0/XI13/MM3_g
+ N_VDD_XI45/XI0/XI13/MM3_s N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI13/MM2 N_XI45/NET277_XI45/XI0/XI13/MM2_d N_NET95_XI45/XI0/XI13/MM2_g
+ N_VDD_XI45/XI0/XI13/MM2_s N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI13/MM1 N_XI45/NET277_XI45/XI0/XI13/MM1_d
+ N_XI45/XI0/NET92_XI45/XI0/XI13/MM1_g N_VDD_XI45/XI0/XI13/MM1_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07
+ PS=5.4e-07
mXI45/XI0/XI13/MM0 N_XI45/NET277_XI45/XI0/XI13/MM0_d
+ N_NET100_XI45/XI0/XI13/MM0_g N_VDD_XI45/XI0/XI13/MM0_s N_VDD_XI10/MM0_b P_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI12/MM3 N_XI45/NET278_XI45/XI0/XI12/MM3_d N_NET79_XI45/XI0/XI12/MM3_g
+ N_VDD_XI45/XI0/XI12/MM3_s N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI12/MM2 N_XI45/NET278_XI45/XI0/XI12/MM2_d
+ N_XI45/XI0/NET081_XI45/XI0/XI12/MM2_g N_VDD_XI45/XI0/XI12/MM2_s
+ N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07
+ PS=5.4e-07
mXI45/XI0/XI12/MM1 N_XI45/NET278_XI45/XI0/XI12/MM1_d
+ N_NET105_XI45/XI0/XI12/MM1_g N_VDD_XI45/XI0/XI12/MM1_s N_VDD_XI10/MM0_b P_18
+ L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI12/MM0 N_XI45/NET278_XI45/XI0/XI12/MM0_d
+ N_NET100_XI45/XI0/XI12/MM0_g N_VDD_XI45/XI0/XI12/MM0_s N_VDD_XI10/MM0_b P_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI11/MM3 N_XI45/NET266_XI45/XI0/XI11/MM3_d N_NET79_XI45/XI0/XI11/MM3_g
+ N_VDD_XI45/XI0/XI11/MM3_s N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI0/XI11/MM2 N_XI45/NET266_XI45/XI0/XI11/MM2_d N_NET95_XI45/XI0/XI11/MM2_g
+ N_VDD_XI45/XI0/XI11/MM2_s N_VDD_XI10/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI11/MM1 N_XI45/NET266_XI45/XI0/XI11/MM1_d
+ N_NET105_XI45/XI0/XI11/MM1_g N_VDD_XI45/XI0/XI11/MM1_s N_VDD_XI10/MM0_b P_18
+ L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI0/XI11/MM0 N_XI45/NET266_XI45/XI0/XI11/MM0_d
+ N_NET100_XI45/XI0/XI11/MM0_g N_VDD_XI45/XI0/XI11/MM0_s N_VDD_XI10/MM0_b P_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI11/MM0 N_XI45/NET252_XI45/XI1/XI11/MM0_d
+ N_NET110_XI45/XI1/XI11/MM0_g N_VDD_XI45/XI1/XI11/MM0_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13
+ PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI11/MM1 N_XI45/NET252_XI45/XI1/XI11/MM1_d N_NET90_XI45/XI1/XI11/MM1_g
+ N_VDD_XI45/XI1/XI11/MM1_s N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI11/MM2 N_XI45/NET252_XI45/XI1/XI11/MM2_d
+ N_NET115_XI45/XI1/XI11/MM2_g N_VDD_XI45/XI1/XI11/MM2_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI11/MM3 N_XI45/NET252_XI45/XI1/XI11/MM3_d N_NET79_XI45/XI1/XI11/MM3_g
+ N_VDD_XI45/XI1/XI11/MM3_s N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI12/MM0 N_XI45/NET264_XI45/XI1/XI12/MM0_d
+ N_NET110_XI45/XI1/XI12/MM0_g N_VDD_XI45/XI1/XI12/MM0_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13
+ PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI12/MM1 N_XI45/NET264_XI45/XI1/XI12/MM1_d N_NET90_XI45/XI1/XI12/MM1_g
+ N_VDD_XI45/XI1/XI12/MM1_s N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI12/MM2 N_XI45/NET264_XI45/XI1/XI12/MM2_d
+ N_XI45/XI1/NET081_XI45/XI1/XI12/MM2_g N_VDD_XI45/XI1/XI12/MM2_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI12/MM3 N_XI45/NET264_XI45/XI1/XI12/MM3_d N_NET79_XI45/XI1/XI12/MM3_g
+ N_VDD_XI45/XI1/XI12/MM3_s N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI13/MM0 N_XI45/NET263_XI45/XI1/XI13/MM0_d
+ N_NET110_XI45/XI1/XI13/MM0_g N_VDD_XI45/XI1/XI13/MM0_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13
+ PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI13/MM1 N_XI45/NET263_XI45/XI1/XI13/MM1_d
+ N_XI45/XI1/NET92_XI45/XI1/XI13/MM1_g N_VDD_XI45/XI1/XI13/MM1_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI13/MM2 N_XI45/NET263_XI45/XI1/XI13/MM2_d
+ N_NET115_XI45/XI1/XI13/MM2_g N_VDD_XI45/XI1/XI13/MM2_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI13/MM3 N_XI45/NET263_XI45/XI1/XI13/MM3_d N_NET79_XI45/XI1/XI13/MM3_g
+ N_VDD_XI45/XI1/XI13/MM3_s N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI14/MM0 N_XI45/NET262_XI45/XI1/XI14/MM0_d
+ N_NET110_XI45/XI1/XI14/MM0_g N_VDD_XI45/XI1/XI14/MM0_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13
+ PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI14/MM1 N_XI45/NET262_XI45/XI1/XI14/MM1_d
+ N_XI45/XI1/NET92_XI45/XI1/XI14/MM1_g N_VDD_XI45/XI1/XI14/MM1_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI14/MM2 N_XI45/NET262_XI45/XI1/XI14/MM2_d
+ N_XI45/XI1/NET081_XI45/XI1/XI14/MM2_g N_VDD_XI45/XI1/XI14/MM2_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI14/MM3 N_XI45/NET262_XI45/XI1/XI14/MM3_d N_NET79_XI45/XI1/XI14/MM3_g
+ N_VDD_XI45/XI1/XI14/MM3_s N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI15/MM0 N_XI45/NET261_XI45/XI1/XI15/MM0_d
+ N_XI45/XI1/NET96_XI45/XI1/XI15/MM0_g N_VDD_XI45/XI1/XI15/MM0_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13
+ PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI15/MM1 N_XI45/NET261_XI45/XI1/XI15/MM1_d N_NET90_XI45/XI1/XI15/MM1_g
+ N_VDD_XI45/XI1/XI15/MM1_s N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI15/MM2 N_XI45/NET261_XI45/XI1/XI15/MM2_d
+ N_NET115_XI45/XI1/XI15/MM2_g N_VDD_XI45/XI1/XI15/MM2_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI15/MM3 N_XI45/NET261_XI45/XI1/XI15/MM3_d N_NET79_XI45/XI1/XI15/MM3_g
+ N_VDD_XI45/XI1/XI15/MM3_s N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI16/MM0 N_XI45/NET260_XI45/XI1/XI16/MM0_d
+ N_XI45/XI1/NET96_XI45/XI1/XI16/MM0_g N_VDD_XI45/XI1/XI16/MM0_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13
+ PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI16/MM1 N_XI45/NET260_XI45/XI1/XI16/MM1_d N_NET90_XI45/XI1/XI16/MM1_g
+ N_VDD_XI45/XI1/XI16/MM1_s N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.269e-13 AS=1.269e-13 PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI16/MM2 N_XI45/NET260_XI45/XI1/XI16/MM2_d
+ N_XI45/XI1/NET081_XI45/XI1/XI16/MM2_g N_VDD_XI45/XI1/XI16/MM2_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI16/MM3 N_XI45/NET260_XI45/XI1/XI16/MM3_d N_NET79_XI45/XI1/XI16/MM3_g
+ N_VDD_XI45/XI1/XI16/MM3_s N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI17/MM0 N_XI45/NET259_XI45/XI1/XI17/MM0_d
+ N_XI45/XI1/NET96_XI45/XI1/XI17/MM0_g N_VDD_XI45/XI1/XI17/MM0_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13
+ PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI17/MM1 N_XI45/NET259_XI45/XI1/XI17/MM1_d
+ N_XI45/XI1/NET92_XI45/XI1/XI17/MM1_g N_VDD_XI45/XI1/XI17/MM1_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI17/MM2 N_XI45/NET259_XI45/XI1/XI17/MM2_d
+ N_NET115_XI45/XI1/XI17/MM2_g N_VDD_XI45/XI1/XI17/MM2_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI17/MM3 N_XI45/NET259_XI45/XI1/XI17/MM3_d N_NET79_XI45/XI1/XI17/MM3_g
+ N_VDD_XI45/XI1/XI17/MM3_s N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI18/MM0 N_XI45/NET258_XI45/XI1/XI18/MM0_d
+ N_XI45/XI1/NET96_XI45/XI1/XI18/MM0_g N_VDD_XI45/XI1/XI18/MM0_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.269e-13
+ PD=1.45e-06 PS=5.4e-07
mXI45/XI1/XI18/MM1 N_XI45/NET258_XI45/XI1/XI18/MM1_d
+ N_XI45/XI1/NET92_XI45/XI1/XI18/MM1_g N_VDD_XI45/XI1/XI18/MM1_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI18/MM2 N_XI45/NET258_XI45/XI1/XI18/MM2_d
+ N_XI45/XI1/NET081_XI45/XI1/XI18/MM2_g N_VDD_XI45/XI1/XI18/MM2_s
+ N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.269e-13
+ PD=5.4e-07 PS=5.4e-07
mXI45/XI1/XI18/MM3 N_XI45/NET258_XI45/XI1/XI18/MM3_d N_NET79_XI45/XI1/XI18/MM3_g
+ N_VDD_XI45/XI1/XI18/MM3_s N_VDD_XI45/XI1/XI11/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
mXI19/MM19 N_XI19/NET37_XI19/MM19_d N_XI19/NET0139_XI19/MM19_g N_VDD_XI19/MM19_s
+ N_VDD_XI19/MM19_b P_18 L=8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI19/XI0/MM0 N_NET79_XI19/XI0/MM0_d N_XI19/NET37_XI19/XI0/MM0_g
+ N_VDD_XI19/XI0/MM0_s N_VDD_XI19/MM19_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=5.325e-13 PD=2.48e-06 PS=7.1e-07
mXI19/XI0/MM1 N_NET79_XI19/XI0/MM1_d N_NET81_XI19/XI0/MM1_g N_VDD_XI19/XI0/MM1_s
+ N_VDD_XI19/MM19_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=5.325e-13
+ PD=2.48e-06 PS=7.1e-07
mXI19/MM24 N_XI19/NET082_XI19/MM24_d N_NET81_XI19/MM24_g N_VDD_XI19/MM24_s
+ N_VDD_XI19/MM19_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI19/MM23 N_XI19/NET086_XI19/MM23_d N_XI19/NET082_XI19/MM23_g N_VDD_XI19/MM23_s
+ N_VDD_XI19/MM19_b P_18 L=3e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI19/MM27 N_NET0265_XI19/MM27_d N_XI19/NET0100_XI19/MM27_g N_VDD_XI19/MM27_s
+ N_VDD_XI19/MM19_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI19/MM29 N_XI19/NET0100_XI19/MM29_d N_NET82_XI19/MM29_g N_VDD_XI19/MM29_s
+ N_VDD_XI19/MM19_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=8.85e-13 PD=2.48e-06
+ PS=2.68e-06
mXI19/MM17 N_NET82_XI19/MM17_d N_XI19/NET9_XI19/MM17_g N_VDD_XI19/MM17_s
+ N_VDD_XI19/MM19_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI19/XI1/MM1 N_XI19/NET9_XI19/XI1/MM1_d N_XI19/NET086_XI19/XI1/MM1_g
+ N_VDD_XI19/XI1/MM1_s N_VDD_XI19/MM19_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=5.325e-13 PD=2.48e-06 PS=7.1e-07
mXI19/XI1/MM0 N_XI19/NET9_XI19/XI1/MM0_d N_XI19/NET086_XI19/XI1/MM0_g
+ N_VDD_XI19/XI1/MM0_s N_VDD_XI19/MM19_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=5.325e-13 PD=2.48e-06 PS=7.1e-07
mXI49/MM1 N_NET0208_XI49/MM1_d N_NET0207_XI49/MM1_g N_VDD_XI49/MM1_s
+ N_VDD_XI49/MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI48/MM1 N_NET0207_XI48/MM1_d N_NET141_XI48/MM1_g N_VDD_XI48/MM1_s
+ N_VDD_XI49/MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI45/XI58/MM3 N_XI45/XI58/NET13_XI45/XI58/MM3_d N_XI45/NET258_XI45/XI58/MM3_g
+ N_VDD_XI45/XI58/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI59/MM3 N_XI45/XI59/NET13_XI45/XI59/MM3_d N_XI45/NET259_XI45/XI59/MM3_g
+ N_VDD_XI45/XI59/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI60/MM3 N_XI45/XI60/NET13_XI45/XI60/MM3_d N_XI45/NET260_XI45/XI60/MM3_g
+ N_VDD_XI45/XI60/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI61/MM3 N_XI45/XI61/NET13_XI45/XI61/MM3_d N_XI45/NET261_XI45/XI61/MM3_g
+ N_VDD_XI45/XI61/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI62/MM3 N_XI45/XI62/NET13_XI45/XI62/MM3_d N_XI45/NET262_XI45/XI62/MM3_g
+ N_VDD_XI45/XI62/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI63/MM3 N_XI45/XI63/NET13_XI45/XI63/MM3_d N_XI45/NET263_XI45/XI63/MM3_g
+ N_VDD_XI45/XI63/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI64/MM3 N_XI45/XI64/NET13_XI45/XI64/MM3_d N_XI45/NET264_XI45/XI64/MM3_g
+ N_VDD_XI45/XI64/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI65/MM3 N_XI45/XI65/NET13_XI45/XI65/MM3_d N_XI45/NET252_XI45/XI65/MM3_g
+ N_VDD_XI45/XI65/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI57/MM3 N_XI45/XI57/NET13_XI45/XI57/MM3_d N_XI45/NET258_XI45/XI57/MM3_g
+ N_VDD_XI45/XI57/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI56/MM3 N_XI45/XI56/NET13_XI45/XI56/MM3_d N_XI45/NET259_XI45/XI56/MM3_g
+ N_VDD_XI45/XI56/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI55/MM3 N_XI45/XI55/NET13_XI45/XI55/MM3_d N_XI45/NET260_XI45/XI55/MM3_g
+ N_VDD_XI45/XI55/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI54/MM3 N_XI45/XI54/NET13_XI45/XI54/MM3_d N_XI45/NET261_XI45/XI54/MM3_g
+ N_VDD_XI45/XI54/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI53/MM3 N_XI45/XI53/NET13_XI45/XI53/MM3_d N_XI45/NET262_XI45/XI53/MM3_g
+ N_VDD_XI45/XI53/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI52/MM3 N_XI45/XI52/NET13_XI45/XI52/MM3_d N_XI45/NET263_XI45/XI52/MM3_g
+ N_VDD_XI45/XI52/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI51/MM3 N_XI45/XI51/NET13_XI45/XI51/MM3_d N_XI45/NET264_XI45/XI51/MM3_g
+ N_VDD_XI45/XI51/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI50/MM3 N_XI45/XI50/NET13_XI45/XI50/MM3_d N_XI45/NET252_XI45/XI50/MM3_g
+ N_VDD_XI45/XI50/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI42/MM3 N_XI45/XI42/NET13_XI45/XI42/MM3_d N_XI45/NET258_XI45/XI42/MM3_g
+ N_VDD_XI45/XI42/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI43/MM3 N_XI45/XI43/NET13_XI45/XI43/MM3_d N_XI45/NET259_XI45/XI43/MM3_g
+ N_VDD_XI45/XI43/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI44/MM3 N_XI45/XI44/NET13_XI45/XI44/MM3_d N_XI45/NET260_XI45/XI44/MM3_g
+ N_VDD_XI45/XI44/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI45/MM3 N_XI45/XI45/NET13_XI45/XI45/MM3_d N_XI45/NET261_XI45/XI45/MM3_g
+ N_VDD_XI45/XI45/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI46/MM3 N_XI45/XI46/NET13_XI45/XI46/MM3_d N_XI45/NET262_XI45/XI46/MM3_g
+ N_VDD_XI45/XI46/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI47/MM3 N_XI45/XI47/NET13_XI45/XI47/MM3_d N_XI45/NET263_XI45/XI47/MM3_g
+ N_VDD_XI45/XI47/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI48/MM3 N_XI45/XI48/NET13_XI45/XI48/MM3_d N_XI45/NET264_XI45/XI48/MM3_g
+ N_VDD_XI45/XI48/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI49/MM3 N_XI45/XI49/NET13_XI45/XI49/MM3_d N_XI45/NET252_XI45/XI49/MM3_g
+ N_VDD_XI45/XI49/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI41/MM3 N_XI45/XI41/NET13_XI45/XI41/MM3_d N_XI45/NET258_XI45/XI41/MM3_g
+ N_VDD_XI45/XI41/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI40/MM3 N_XI45/XI40/NET13_XI45/XI40/MM3_d N_XI45/NET259_XI45/XI40/MM3_g
+ N_VDD_XI45/XI40/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI39/MM3 N_XI45/XI39/NET13_XI45/XI39/MM3_d N_XI45/NET260_XI45/XI39/MM3_g
+ N_VDD_XI45/XI39/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI38/MM3 N_XI45/XI38/NET13_XI45/XI38/MM3_d N_XI45/NET261_XI45/XI38/MM3_g
+ N_VDD_XI45/XI38/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI37/MM3 N_XI45/XI37/NET13_XI45/XI37/MM3_d N_XI45/NET262_XI45/XI37/MM3_g
+ N_VDD_XI45/XI37/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI36/MM3 N_XI45/XI36/NET13_XI45/XI36/MM3_d N_XI45/NET263_XI45/XI36/MM3_g
+ N_VDD_XI45/XI36/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI35/MM3 N_XI45/XI35/NET13_XI45/XI35/MM3_d N_XI45/NET264_XI45/XI35/MM3_g
+ N_VDD_XI45/XI35/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI34/MM3 N_XI45/XI34/NET13_XI45/XI34/MM3_d N_XI45/NET252_XI45/XI34/MM3_g
+ N_VDD_XI45/XI34/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI26/MM3 N_XI45/XI26/NET13_XI45/XI26/MM3_d N_XI45/NET258_XI45/XI26/MM3_g
+ N_VDD_XI45/XI26/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI27/MM3 N_XI45/XI27/NET13_XI45/XI27/MM3_d N_XI45/NET259_XI45/XI27/MM3_g
+ N_VDD_XI45/XI27/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI28/MM3 N_XI45/XI28/NET13_XI45/XI28/MM3_d N_XI45/NET260_XI45/XI28/MM3_g
+ N_VDD_XI45/XI28/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI29/MM3 N_XI45/XI29/NET13_XI45/XI29/MM3_d N_XI45/NET261_XI45/XI29/MM3_g
+ N_VDD_XI45/XI29/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI30/MM3 N_XI45/XI30/NET13_XI45/XI30/MM3_d N_XI45/NET262_XI45/XI30/MM3_g
+ N_VDD_XI45/XI30/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI31/MM3 N_XI45/XI31/NET13_XI45/XI31/MM3_d N_XI45/NET263_XI45/XI31/MM3_g
+ N_VDD_XI45/XI31/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI32/MM3 N_XI45/XI32/NET13_XI45/XI32/MM3_d N_XI45/NET264_XI45/XI32/MM3_g
+ N_VDD_XI45/XI32/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI33/MM3 N_XI45/XI33/NET13_XI45/XI33/MM3_d N_XI45/NET252_XI45/XI33/MM3_g
+ N_VDD_XI45/XI33/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI25/MM3 N_XI45/XI25/NET13_XI45/XI25/MM3_d N_XI45/NET258_XI45/XI25/MM3_g
+ N_VDD_XI45/XI25/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI24/MM3 N_XI45/XI24/NET13_XI45/XI24/MM3_d N_XI45/NET259_XI45/XI24/MM3_g
+ N_VDD_XI45/XI24/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI23/MM3 N_XI45/XI23/NET13_XI45/XI23/MM3_d N_XI45/NET260_XI45/XI23/MM3_g
+ N_VDD_XI45/XI23/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI22/MM3 N_XI45/XI22/NET13_XI45/XI22/MM3_d N_XI45/NET261_XI45/XI22/MM3_g
+ N_VDD_XI45/XI22/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI21/MM3 N_XI45/XI21/NET13_XI45/XI21/MM3_d N_XI45/NET262_XI45/XI21/MM3_g
+ N_VDD_XI45/XI21/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI20/MM3 N_XI45/XI20/NET13_XI45/XI20/MM3_d N_XI45/NET263_XI45/XI20/MM3_g
+ N_VDD_XI45/XI20/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI19/MM3 N_XI45/XI19/NET13_XI45/XI19/MM3_d N_XI45/NET264_XI45/XI19/MM3_g
+ N_VDD_XI45/XI19/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI18/MM3 N_XI45/XI18/NET13_XI45/XI18/MM3_d N_XI45/NET252_XI45/XI18/MM3_g
+ N_VDD_XI45/XI18/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI10/MM3 N_XI45/XI10/NET13_XI45/XI10/MM3_d N_XI45/NET258_XI45/XI10/MM3_g
+ N_VDD_XI45/XI10/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI11/MM3 N_XI45/XI11/NET13_XI45/XI11/MM3_d N_XI45/NET259_XI45/XI11/MM3_g
+ N_VDD_XI45/XI11/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI12/MM3 N_XI45/XI12/NET13_XI45/XI12/MM3_d N_XI45/NET260_XI45/XI12/MM3_g
+ N_VDD_XI45/XI12/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI13/MM3 N_XI45/XI13/NET13_XI45/XI13/MM3_d N_XI45/NET261_XI45/XI13/MM3_g
+ N_VDD_XI45/XI13/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI14/MM3 N_XI45/XI14/NET13_XI45/XI14/MM3_d N_XI45/NET262_XI45/XI14/MM3_g
+ N_VDD_XI45/XI14/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI15/MM3 N_XI45/XI15/NET13_XI45/XI15/MM3_d N_XI45/NET263_XI45/XI15/MM3_g
+ N_VDD_XI45/XI15/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI16/MM3 N_XI45/XI16/NET13_XI45/XI16/MM3_d N_XI45/NET264_XI45/XI16/MM3_g
+ N_VDD_XI45/XI16/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI17/MM3 N_XI45/XI17/NET13_XI45/XI17/MM3_d N_XI45/NET252_XI45/XI17/MM3_g
+ N_VDD_XI45/XI17/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI9/MM3 N_XI45/XI9/NET13_XI45/XI9/MM3_d N_XI45/NET258_XI45/XI9/MM3_g
+ N_VDD_XI45/XI9/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI8/MM3 N_XI45/XI8/NET13_XI45/XI8/MM3_d N_XI45/NET259_XI45/XI8/MM3_g
+ N_VDD_XI45/XI8/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI7/MM3 N_XI45/XI7/NET13_XI45/XI7/MM3_d N_XI45/NET260_XI45/XI7/MM3_g
+ N_VDD_XI45/XI7/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI6/MM3 N_XI45/XI6/NET13_XI45/XI6/MM3_d N_XI45/NET261_XI45/XI6/MM3_g
+ N_VDD_XI45/XI6/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI5/MM3 N_XI45/XI5/NET13_XI45/XI5/MM3_d N_XI45/NET262_XI45/XI5/MM3_g
+ N_VDD_XI45/XI5/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI4/MM3 N_XI45/XI4/NET13_XI45/XI4/MM3_d N_XI45/NET263_XI45/XI4/MM3_g
+ N_VDD_XI45/XI4/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI3/MM3 N_XI45/XI3/NET13_XI45/XI3/MM3_d N_XI45/NET264_XI45/XI3/MM3_g
+ N_VDD_XI45/XI3/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI2/MM3 N_XI45/XI2/NET13_XI45/XI2/MM3_d N_XI45/NET252_XI45/XI2/MM3_g
+ N_VDD_XI45/XI2/MM3_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.303e-13 PD=7.2e-07 PS=1.45e-06
mXI45/XI58/MM2 N_NET10_XI45/XI58/MM2_d N_XI45/NET272_XI45/XI58/MM2_g
+ N_XI45/XI58/NET13_XI45/XI58/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI59/MM2 N_NET11_XI45/XI59/MM2_d N_XI45/NET272_XI45/XI59/MM2_g
+ N_XI45/XI59/NET13_XI45/XI59/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI60/MM2 N_NET12_XI45/XI60/MM2_d N_XI45/NET272_XI45/XI60/MM2_g
+ N_XI45/XI60/NET13_XI45/XI60/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI61/MM2 N_NET13_XI45/XI61/MM2_d N_XI45/NET272_XI45/XI61/MM2_g
+ N_XI45/XI61/NET13_XI45/XI61/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI62/MM2 N_NET14_XI45/XI62/MM2_d N_XI45/NET272_XI45/XI62/MM2_g
+ N_XI45/XI62/NET13_XI45/XI62/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI63/MM2 N_NET15_XI45/XI63/MM2_d N_XI45/NET272_XI45/XI63/MM2_g
+ N_XI45/XI63/NET13_XI45/XI63/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI64/MM2 N_NET16_XI45/XI64/MM2_d N_XI45/NET272_XI45/XI64/MM2_g
+ N_XI45/XI64/NET13_XI45/XI64/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI65/MM2 N_NET17_XI45/XI65/MM2_d N_XI45/NET272_XI45/XI65/MM2_g
+ N_XI45/XI65/NET13_XI45/XI65/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI57/MM2 N_NET18_XI45/XI57/MM2_d N_XI45/NET273_XI45/XI57/MM2_g
+ N_XI45/XI57/NET13_XI45/XI57/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI56/MM2 N_NET19_XI45/XI56/MM2_d N_XI45/NET273_XI45/XI56/MM2_g
+ N_XI45/XI56/NET13_XI45/XI56/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI55/MM2 N_NET20_XI45/XI55/MM2_d N_XI45/NET273_XI45/XI55/MM2_g
+ N_XI45/XI55/NET13_XI45/XI55/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI54/MM2 N_NET21_XI45/XI54/MM2_d N_XI45/NET273_XI45/XI54/MM2_g
+ N_XI45/XI54/NET13_XI45/XI54/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI53/MM2 N_NET22_XI45/XI53/MM2_d N_XI45/NET273_XI45/XI53/MM2_g
+ N_XI45/XI53/NET13_XI45/XI53/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI52/MM2 N_NET23_XI45/XI52/MM2_d N_XI45/NET273_XI45/XI52/MM2_g
+ N_XI45/XI52/NET13_XI45/XI52/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI51/MM2 N_NET24_XI45/XI51/MM2_d N_XI45/NET273_XI45/XI51/MM2_g
+ N_XI45/XI51/NET13_XI45/XI51/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI50/MM2 N_NET25_XI45/XI50/MM2_d N_XI45/NET273_XI45/XI50/MM2_g
+ N_XI45/XI50/NET13_XI45/XI50/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI42/MM2 N_NET26_XI45/XI42/MM2_d N_XI45/NET274_XI45/XI42/MM2_g
+ N_XI45/XI42/NET13_XI45/XI42/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI43/MM2 N_NET27_XI45/XI43/MM2_d N_XI45/NET274_XI45/XI43/MM2_g
+ N_XI45/XI43/NET13_XI45/XI43/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI44/MM2 N_NET28_XI45/XI44/MM2_d N_XI45/NET274_XI45/XI44/MM2_g
+ N_XI45/XI44/NET13_XI45/XI44/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI45/MM2 N_NET29_XI45/XI45/MM2_d N_XI45/NET274_XI45/XI45/MM2_g
+ N_XI45/XI45/NET13_XI45/XI45/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI46/MM2 N_NET30_XI45/XI46/MM2_d N_XI45/NET274_XI45/XI46/MM2_g
+ N_XI45/XI46/NET13_XI45/XI46/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI47/MM2 N_NET31_XI45/XI47/MM2_d N_XI45/NET274_XI45/XI47/MM2_g
+ N_XI45/XI47/NET13_XI45/XI47/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI48/MM2 N_NET32_XI45/XI48/MM2_d N_XI45/NET274_XI45/XI48/MM2_g
+ N_XI45/XI48/NET13_XI45/XI48/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI49/MM2 N_NET33_XI45/XI49/MM2_d N_XI45/NET274_XI45/XI49/MM2_g
+ N_XI45/XI49/NET13_XI45/XI49/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI41/MM2 N_NET34_XI45/XI41/MM2_d N_XI45/NET275_XI45/XI41/MM2_g
+ N_XI45/XI41/NET13_XI45/XI41/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI40/MM2 N_NET35_XI45/XI40/MM2_d N_XI45/NET275_XI45/XI40/MM2_g
+ N_XI45/XI40/NET13_XI45/XI40/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI39/MM2 N_NET36_XI45/XI39/MM2_d N_XI45/NET275_XI45/XI39/MM2_g
+ N_XI45/XI39/NET13_XI45/XI39/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI38/MM2 N_NET37_XI45/XI38/MM2_d N_XI45/NET275_XI45/XI38/MM2_g
+ N_XI45/XI38/NET13_XI45/XI38/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI37/MM2 N_NET38_XI45/XI37/MM2_d N_XI45/NET275_XI45/XI37/MM2_g
+ N_XI45/XI37/NET13_XI45/XI37/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI36/MM2 N_NET39_XI45/XI36/MM2_d N_XI45/NET275_XI45/XI36/MM2_g
+ N_XI45/XI36/NET13_XI45/XI36/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI35/MM2 N_NET40_XI45/XI35/MM2_d N_XI45/NET275_XI45/XI35/MM2_g
+ N_XI45/XI35/NET13_XI45/XI35/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI34/MM2 N_NET41_XI45/XI34/MM2_d N_XI45/NET275_XI45/XI34/MM2_g
+ N_XI45/XI34/NET13_XI45/XI34/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI26/MM2 N_NET42_XI45/XI26/MM2_d N_XI45/NET276_XI45/XI26/MM2_g
+ N_XI45/XI26/NET13_XI45/XI26/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI27/MM2 N_NET43_XI45/XI27/MM2_d N_XI45/NET276_XI45/XI27/MM2_g
+ N_XI45/XI27/NET13_XI45/XI27/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI28/MM2 N_NET44_XI45/XI28/MM2_d N_XI45/NET276_XI45/XI28/MM2_g
+ N_XI45/XI28/NET13_XI45/XI28/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI29/MM2 N_NET45_XI45/XI29/MM2_d N_XI45/NET276_XI45/XI29/MM2_g
+ N_XI45/XI29/NET13_XI45/XI29/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI30/MM2 N_NET46_XI45/XI30/MM2_d N_XI45/NET276_XI45/XI30/MM2_g
+ N_XI45/XI30/NET13_XI45/XI30/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI31/MM2 N_NET47_XI45/XI31/MM2_d N_XI45/NET276_XI45/XI31/MM2_g
+ N_XI45/XI31/NET13_XI45/XI31/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI32/MM2 N_NET48_XI45/XI32/MM2_d N_XI45/NET276_XI45/XI32/MM2_g
+ N_XI45/XI32/NET13_XI45/XI32/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI33/MM2 N_NET49_XI45/XI33/MM2_d N_XI45/NET276_XI45/XI33/MM2_g
+ N_XI45/XI33/NET13_XI45/XI33/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI25/MM2 N_NET50_XI45/XI25/MM2_d N_XI45/NET277_XI45/XI25/MM2_g
+ N_XI45/XI25/NET13_XI45/XI25/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI24/MM2 N_NET51_XI45/XI24/MM2_d N_XI45/NET277_XI45/XI24/MM2_g
+ N_XI45/XI24/NET13_XI45/XI24/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI23/MM2 N_NET52_XI45/XI23/MM2_d N_XI45/NET277_XI45/XI23/MM2_g
+ N_XI45/XI23/NET13_XI45/XI23/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI22/MM2 N_NET53_XI45/XI22/MM2_d N_XI45/NET277_XI45/XI22/MM2_g
+ N_XI45/XI22/NET13_XI45/XI22/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI21/MM2 N_NET54_XI45/XI21/MM2_d N_XI45/NET277_XI45/XI21/MM2_g
+ N_XI45/XI21/NET13_XI45/XI21/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI20/MM2 N_NET55_XI45/XI20/MM2_d N_XI45/NET277_XI45/XI20/MM2_g
+ N_XI45/XI20/NET13_XI45/XI20/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI19/MM2 N_NET56_XI45/XI19/MM2_d N_XI45/NET277_XI45/XI19/MM2_g
+ N_XI45/XI19/NET13_XI45/XI19/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI18/MM2 N_NET57_XI45/XI18/MM2_d N_XI45/NET277_XI45/XI18/MM2_g
+ N_XI45/XI18/NET13_XI45/XI18/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI10/MM2 N_NET58_XI45/XI10/MM2_d N_XI45/NET278_XI45/XI10/MM2_g
+ N_XI45/XI10/NET13_XI45/XI10/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI11/MM2 N_NET59_XI45/XI11/MM2_d N_XI45/NET278_XI45/XI11/MM2_g
+ N_XI45/XI11/NET13_XI45/XI11/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI12/MM2 N_NET60_XI45/XI12/MM2_d N_XI45/NET278_XI45/XI12/MM2_g
+ N_XI45/XI12/NET13_XI45/XI12/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI13/MM2 N_NET61_XI45/XI13/MM2_d N_XI45/NET278_XI45/XI13/MM2_g
+ N_XI45/XI13/NET13_XI45/XI13/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI14/MM2 N_NET62_XI45/XI14/MM2_d N_XI45/NET278_XI45/XI14/MM2_g
+ N_XI45/XI14/NET13_XI45/XI14/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI15/MM2 N_NET63_XI45/XI15/MM2_d N_XI45/NET278_XI45/XI15/MM2_g
+ N_XI45/XI15/NET13_XI45/XI15/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI16/MM2 N_NET64_XI45/XI16/MM2_d N_XI45/NET278_XI45/XI16/MM2_g
+ N_XI45/XI16/NET13_XI45/XI16/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI17/MM2 N_NET65_XI45/XI17/MM2_d N_XI45/NET278_XI45/XI17/MM2_g
+ N_XI45/XI17/NET13_XI45/XI17/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI9/MM2 N_NET66_XI45/XI9/MM2_d N_XI45/NET266_XI45/XI9/MM2_g
+ N_XI45/XI9/NET13_XI45/XI9/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI8/MM2 N_NET67_XI45/XI8/MM2_d N_XI45/NET266_XI45/XI8/MM2_g
+ N_XI45/XI8/NET13_XI45/XI8/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI7/MM2 N_NET68_XI45/XI7/MM2_d N_XI45/NET266_XI45/XI7/MM2_g
+ N_XI45/XI7/NET13_XI45/XI7/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI6/MM2 N_NET69_XI45/XI6/MM2_d N_XI45/NET266_XI45/XI6/MM2_g
+ N_XI45/XI6/NET13_XI45/XI6/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI5/MM2 N_NET70_XI45/XI5/MM2_d N_XI45/NET266_XI45/XI5/MM2_g
+ N_XI45/XI5/NET13_XI45/XI5/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI4/MM2 N_NET71_XI45/XI4/MM2_d N_XI45/NET266_XI45/XI4/MM2_g
+ N_XI45/XI4/NET13_XI45/XI4/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI3/MM2 N_NET72_XI45/XI3/MM2_d N_XI45/NET266_XI45/XI3/MM2_g
+ N_XI45/XI3/NET13_XI45/XI3/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI45/XI2/MM2 N_NET8_XI45/XI2/MM2_d N_XI45/NET266_XI45/XI2/MM2_g
+ N_XI45/XI2/NET13_XI45/XI2/MM2_s N_VDD_XI45/XI58/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.692e-13 PD=1.45e-06 PS=7.2e-07
mXI7/MM5 N_XI7/NET48_XI7/MM5_d N_NET120_XI7/MM5_g N_VDD_XI7/MM5_s
+ N_VDD_XI7/MM5_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI7/MM7 N_XI7/NET68_XI7/MM7_d N_NET125_XI7/MM7_g N_VDD_XI7/MM7_s
+ N_VDD_XI7/MM5_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI8/MM6 N_NET141_XI8/MM6_d N_NET0174_XI8/MM6_g N_VDD_XI8/MM6_s N_VDD_XI7/MM5_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.5e-12 AS=1.1775e-12 PD=4e-06 PS=2.385e-06
mXI8/MM7 N_NET0174_XI8/MM7_d N_NET141_XI8/MM7_g N_VDD_XI8/MM7_s N_VDD_XI7/MM5_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.27875e-12 PD=3.98e-06 PS=2.4525e-06
mXI7/MM8 N_XI7/NET76_XI7/MM8_d N_NET85_XI7/MM8_g N_VDD_XI7/MM8_s N_VDD_XI7/MM5_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI7/MM0 N_XI7/NET141_XI7/MM0_d N_XI7/NET48_XI7/MM0_g N_NET147_XI7/MM0_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI6/MM0 N_NET147_XI6/MM0_d N_NET81_XI6/MM0_g N_VDD_XI6/MM0_s N_VDD_XI7/MM0_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI8/MM5 N_NET141_XI8/MM5_d N_NET82_XI8/MM5_g N_VDD_XI8/MM5_s N_VDD_XI7/MM5_b
+ P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=3.925e-13 PD=1.98e-06 PS=7.95e-07
mXI8/MM8 N_NET0174_XI8/MM8_d N_NET82_XI8/MM8_g N_VDD_XI8/MM8_s N_VDD_XI7/MM5_b
+ P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.2625e-13 PD=1.98e-06 PS=8.175e-07
mXI7/MM3 N_XI7/NET141_XI7/MM3_d N_NET120_XI7/MM3_g N_NET148_XI7/MM3_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI6/MM1 N_NET148_XI6/MM1_d N_NET81_XI6/MM1_g N_VDD_XI6/MM1_s N_VDD_XI7/MM0_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI7/MM25 N_XI7/NET101_XI7/MM25_d N_XI7/NET68_XI7/MM25_g N_XI7/NET141_XI7/MM25_s
+ N_VDD_XI7/MM25_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI7/MM24 N_XI7/NET101_XI7/MM24_d N_NET125_XI7/MM24_g N_XI7/NET125_XI7/MM24_s
+ N_VDD_XI7/MM25_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI7/MM13 N_XI7/NET125_XI7/MM13_d N_XI7/NET48_XI7/MM13_g N_NET149_XI7/MM13_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI6/MM2 N_NET149_XI6/MM2_d N_NET81_XI6/MM2_g N_VDD_XI6/MM2_s N_VDD_XI7/MM0_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI7/MM12 N_XI7/NET125_XI7/MM12_d N_NET120_XI7/MM12_g N_NET151_XI7/MM12_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI6/MM3 N_NET151_XI6/MM3_d N_NET81_XI6/MM3_g N_VDD_XI6/MM3_s N_VDD_XI7/MM0_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI7/MM32 N_NET139_XI7/MM32_d N_XI7/NET76_XI7/MM32_g N_XI7/NET101_XI7/MM32_s
+ N_VDD_XI7/MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI7/MM33 N_NET139_XI7/MM33_d N_NET85_XI7/MM33_g N_XI7/NET89_XI7/MM33_s
+ N_VDD_XI7/MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI7/MM14 N_XI7/NET113_XI7/MM14_d N_XI7/NET48_XI7/MM14_g N_NET152_XI7/MM14_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI6/MM5 N_NET152_XI6/MM5_d N_NET81_XI6/MM5_g N_VDD_XI6/MM5_s N_VDD_XI7/MM0_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI7/MM15 N_XI7/NET113_XI7/MM15_d N_NET120_XI7/MM15_g N_NET153_XI7/MM15_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI6/MM7 N_NET153_XI6/MM7_d N_NET81_XI6/MM7_g N_VDD_XI6/MM7_s N_VDD_XI7/MM0_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI50/MM1 N_NET0215_XI50/MM1_d N_NET0214_XI50/MM1_g N_VDD_XI50/MM1_s
+ N_VDD_XI7/MM5_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI51/MM1 N_NET0214_XI51/MM1_d N_NET134_XI51/MM1_g N_VDD_XI51/MM1_s
+ N_VDD_XI7/MM5_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI7/MM28 N_XI7/NET89_XI7/MM28_d N_XI7/NET68_XI7/MM28_g N_XI7/NET113_XI7/MM28_s
+ N_VDD_XI7/MM25_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI7/MM29 N_XI7/NET89_XI7/MM29_d N_NET125_XI7/MM29_g N_XI7/NET109_XI7/MM29_s
+ N_VDD_XI7/MM25_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI7/MM21 N_XI7/NET109_XI7/MM21_d N_XI7/NET48_XI7/MM21_g N_NET154_XI7/MM21_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI6/MM6 N_NET154_XI6/MM6_d N_NET81_XI6/MM6_g N_VDD_XI6/MM6_s N_VDD_XI7/MM0_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI7/MM20 N_XI7/NET109_XI7/MM20_d N_NET120_XI7/MM20_g N_NET155_XI7/MM20_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI6/MM4 N_NET155_XI6/MM4_d N_NET81_XI6/MM4_g N_VDD_XI6/MM4_s N_VDD_XI7/MM0_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI7/MM61 N_XI7/NET29_XI7/MM61_d N_XI7/NET48_XI7/MM61_g N_NET156_XI7/MM61_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI6/MM13 N_NET156_XI6/MM13_d N_NET81_XI6/MM13_g N_VDD_XI6/MM13_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM60 N_XI7/NET29_XI7/MM60_d N_NET120_XI7/MM60_g N_NET157_XI7/MM60_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI6/MM15 N_NET157_XI6/MM15_d N_NET81_XI6/MM15_g N_VDD_XI6/MM15_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM52 N_XI7/NET57_XI7/MM52_d N_XI7/NET68_XI7/MM52_g N_XI7/NET29_XI7/MM52_s
+ N_VDD_XI7/MM25_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI7/MM53 N_XI7/NET57_XI7/MM53_d N_NET125_XI7/MM53_g N_XI7/NET33_XI7/MM53_s
+ N_VDD_XI7/MM25_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI7/MM58 N_XI7/NET33_XI7/MM58_d N_XI7/NET48_XI7/MM58_g N_NET150_XI7/MM58_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI6/MM14 N_NET150_XI6/MM14_d N_NET81_XI6/MM14_g N_VDD_XI6/MM14_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM59 N_XI7/NET33_XI7/MM59_d N_NET120_XI7/MM59_g N_NET158_XI7/MM59_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI6/MM12 N_NET158_XI6/MM12_d N_NET81_XI6/MM12_g N_VDD_XI6/MM12_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM49 N_NET165_XI7/MM49_d N_XI7/NET76_XI7/MM49_g N_XI7/NET57_XI7/MM49_s
+ N_VDD_XI7/MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI9/MM6 N_NET134_XI9/MM6_d N_NET0181_XI9/MM6_g N_VDD_XI9/MM6_s N_VDD_XI9/MM6_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.5e-12 AS=1.1775e-12 PD=4e-06 PS=2.385e-06
mXI9/MM7 N_NET0181_XI9/MM7_d N_NET134_XI9/MM7_g N_VDD_XI9/MM7_s N_VDD_XI9/MM6_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.27875e-12 PD=3.98e-06 PS=2.4525e-06
mXI7/MM48 N_NET165_XI7/MM48_d N_NET85_XI7/MM48_g N_XI7/NET69_XI7/MM48_s
+ N_VDD_XI7/MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI7/MM57 N_XI7/NET45_XI7/MM57_d N_XI7/NET48_XI7/MM57_g N_NET159_XI7/MM57_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI6/MM10 N_NET159_XI6/MM10_d N_NET81_XI6/MM10_g N_VDD_XI6/MM10_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI7/MM56 N_XI7/NET45_XI7/MM56_d N_NET120_XI7/MM56_g N_NET160_XI7/MM56_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI6/MM8 N_NET160_XI6/MM8_d N_NET81_XI6/MM8_g N_VDD_XI6/MM8_s N_VDD_XI7/MM0_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI7/MM51 N_XI7/NET69_XI7/MM51_d N_XI7/NET68_XI7/MM51_g N_XI7/NET45_XI7/MM51_s
+ N_VDD_XI7/MM25_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI9/MM5 N_NET134_XI9/MM5_d N_NET82_XI9/MM5_g N_VDD_XI9/MM5_s N_VDD_XI9/MM6_b
+ P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=3.925e-13 PD=1.98e-06 PS=7.95e-07
mXI9/MM8 N_NET0181_XI9/MM8_d N_NET82_XI9/MM8_g N_VDD_XI9/MM8_s N_VDD_XI9/MM6_b
+ P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.2625e-13 PD=1.98e-06 PS=8.175e-07
mXI7/MM50 N_XI7/NET69_XI7/MM50_d N_NET125_XI7/MM50_g N_XI7/NET49_XI7/MM50_s
+ N_VDD_XI7/MM25_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI7/MM54 N_XI7/NET49_XI7/MM54_d N_XI7/NET48_XI7/MM54_g N_NET161_XI7/MM54_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI6/MM9 N_NET161_XI6/MM9_d N_NET81_XI6/MM9_g N_VDD_XI6/MM9_s N_VDD_XI7/MM0_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI7/MM55 N_XI7/NET49_XI7/MM55_d N_NET120_XI7/MM55_g N_NET162_XI7/MM55_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
mXI6/MM11 N_NET162_XI6/MM11_d N_NET81_XI6/MM11_g N_VDD_XI6/MM11_s
+ N_VDD_XI7/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
c_1 XI5/NET02326 0 0.148602f
c_2 XI5/NET02370 0 0.148602f
c_3 XI5/NET02402 0 0.148602f
c_4 XI5/NET02434 0 0.148602f
c_5 XI5/NET02466 0 0.148602f
c_6 XI5/NET04286 0 0.148602f
c_7 XI5/NET04318 0 0.148602f
c_8 XI5/NET03466 0 0.148602f
c_9 XI5/NET05406 0 0.148602f
c_10 XI5/NET05362 0 0.148602f
c_11 XI5/NET05318 0 0.148602f
c_12 XI5/NET05286 0 0.148602f
c_13 XI5/NET05254 0 0.148602f
c_14 XI5/NET05222 0 0.148602f
c_15 XI5/NET05182 0 0.148602f
c_16 XI5/NET05150 0 0.148602f
c_17 XI5/NET05114 0 0.148602f
c_18 XI5/NET05082 0 0.148602f
c_19 XI5/NET05050 0 0.148602f
c_20 XI5/NET05018 0 0.148602f
c_21 XI5/NET04986 0 0.148602f
c_22 XI5/NET04954 0 0.148602f
c_23 XI5/NET04914 0 0.148602f
c_24 XI5/NET04882 0 0.148602f
c_25 XI5/NET04850 0 0.148602f
c_26 XI5/NET04818 0 0.148602f
c_27 XI5/NET04766 0 0.148602f
c_28 XI5/NET04734 0 0.148602f
c_29 XI5/NET04654 0 0.148602f
c_30 XI5/NET04618 0 0.148602f
c_31 XI5/NET04586 0 0.148602f
c_32 XI5/NET04390 0 0.148602f
c_33 XI5/NET01346 0 0.180551f
c_34 XI5/NET01378 0 0.176433f
c_35 XI5/NET01410 0 0.176433f
c_36 XI5/NET01442 0 0.176433f
c_37 XI5/NET01474 0 0.176433f
c_38 XI5/NET01506 0 0.176433f
c_39 XI5/NET01538 0 0.176433f
c_40 XI5/NET01570 0 0.176433f
c_41 XI5/NET01602 0 0.18066f
c_42 XI5/NET01634 0 0.176433f
c_43 XI5/NET01666 0 0.176433f
c_44 XI5/NET01698 0 0.176433f
c_45 XI5/NET01730 0 0.176433f
c_46 XI5/NET01762 0 0.176433f
c_47 XI5/NET01794 0 0.176433f
c_48 XI5/NET01826 0 0.176433f
c_49 XI5/NET01858 0 0.18066f
c_50 XI5/NET01890 0 0.176433f
c_51 XI5/NET01922 0 0.176433f
c_52 XI5/NET01954 0 0.176433f
c_53 XI5/NET01986 0 0.176433f
c_54 XI5/NET02018 0 0.176433f
c_55 XI5/NET02050 0 0.176433f
c_56 XI5/NET02082 0 0.176433f
c_57 XI5/NET02114 0 0.18066f
c_58 XI5/NET02146 0 0.176433f
c_59 XI5/NET02178 0 0.176433f
c_60 XI5/NET02210 0 0.176433f
c_61 XI5/NET02242 0 0.176433f
c_62 XI5/NET02274 0 0.176433f
c_63 XI5/NET02278 0 0.176433f
c_64 XI5/NET04538 0 0.176433f
c_65 XI5/NET02310 0 0.176433f
c_66 XI5/NET02366 0 0.176433f
c_67 XI5/NET02398 0 0.176433f
c_68 XI5/NET02430 0 0.176433f
c_69 XI5/NET02462 0 0.176433f
c_70 XI5/NET04282 0 0.176433f
c_71 XI5/NET04314 0 0.176433f
c_72 XI5/NET03462 0 0.176433f
c_73 XI5/NET05402 0 0.176433f
c_74 XI5/NET05358 0 0.176433f
c_75 XI5/NET05314 0 0.176433f
c_76 XI5/NET05282 0 0.176433f
c_77 XI5/NET05250 0 0.176433f
c_78 XI5/NET05218 0 0.176433f
c_79 XI5/NET05178 0 0.176433f
c_80 XI5/NET05146 0 0.176433f
c_81 XI5/NET05110 0 0.176433f
c_82 XI5/NET05078 0 0.176433f
c_83 XI5/NET05046 0 0.176433f
c_84 XI5/NET05014 0 0.176433f
c_85 XI5/NET04982 0 0.176433f
c_86 XI5/NET04950 0 0.176433f
c_87 XI5/NET04910 0 0.176433f
c_88 XI5/NET04878 0 0.176433f
c_89 XI5/NET04846 0 0.176433f
c_90 XI5/NET04814 0 0.176433f
c_91 XI5/NET04762 0 0.176433f
c_92 XI5/NET04730 0 0.176433f
c_93 XI5/NET04650 0 0.176433f
c_94 XI5/NET04614 0 0.176433f
c_95 XI5/NET04582 0 0.176433f
c_96 XI5/NET04386 0 0.176433f
c_97 XI5/NET01342 0 0.180551f
c_98 XI5/NET01374 0 0.176433f
c_99 XI5/NET01406 0 0.176433f
c_100 XI5/NET01438 0 0.176433f
c_101 XI5/NET01470 0 0.176433f
c_102 XI5/NET01502 0 0.176433f
c_103 XI5/NET01534 0 0.176433f
c_104 XI5/NET01566 0 0.176433f
c_105 XI5/NET01598 0 0.18066f
c_106 XI5/NET01630 0 0.176433f
c_107 XI5/NET01662 0 0.176433f
c_108 XI5/NET01694 0 0.176433f
c_109 XI5/NET01726 0 0.176433f
c_110 XI5/NET01758 0 0.176433f
c_111 XI5/NET01790 0 0.176433f
c_112 XI5/NET01822 0 0.176433f
c_113 XI5/NET01854 0 0.18066f
c_114 XI5/NET01886 0 0.176433f
c_115 XI5/NET01918 0 0.176433f
c_116 XI5/NET01950 0 0.176433f
c_117 XI5/NET01982 0 0.176433f
c_118 XI5/NET02014 0 0.176433f
c_119 XI5/NET02046 0 0.176433f
c_120 XI5/NET02078 0 0.176433f
c_121 XI5/NET02110 0 0.18066f
c_122 XI5/NET02142 0 0.176433f
c_123 XI5/NET02174 0 0.176433f
c_124 XI5/NET02206 0 0.176433f
c_125 XI5/NET02238 0 0.176433f
c_126 XI5/NET02270 0 0.176433f
c_127 XI5/NET02282 0 0.176433f
c_128 XI5/NET04534 0 0.176433f
c_129 XI5/NET02338 0 0.176433f
c_130 XI5/NET02362 0 0.176433f
c_131 XI5/NET02394 0 0.176433f
c_132 XI5/NET02426 0 0.176433f
c_133 XI5/NET02458 0 0.176433f
c_134 XI5/NET04278 0 0.176433f
c_135 XI5/NET04310 0 0.176433f
c_136 XI5/NET03458 0 0.176433f
c_137 XI5/NET05398 0 0.176433f
c_138 XI5/NET05354 0 0.176433f
c_139 XI5/NET05310 0 0.176433f
c_140 XI5/NET05278 0 0.176433f
c_141 XI5/NET05246 0 0.176433f
c_142 XI5/NET05214 0 0.176433f
c_143 XI5/NET05174 0 0.176433f
c_144 XI5/NET05142 0 0.176433f
c_145 XI5/NET05106 0 0.176433f
c_146 XI5/NET05074 0 0.176433f
c_147 XI5/NET05042 0 0.176433f
c_148 XI5/NET05010 0 0.176433f
c_149 XI5/NET04978 0 0.176433f
c_150 XI5/NET04946 0 0.176433f
c_151 XI5/NET04906 0 0.176433f
c_152 XI5/NET04874 0 0.176433f
c_153 XI5/NET04842 0 0.176433f
c_154 XI5/NET04810 0 0.176433f
c_155 XI5/NET04758 0 0.176433f
c_156 XI5/NET04722 0 0.176433f
c_157 XI5/NET04642 0 0.176433f
c_158 XI5/NET04610 0 0.176433f
c_159 XI5/NET04578 0 0.176433f
c_160 XI5/NET04382 0 0.176433f
c_161 XI5/NET01338 0 0.180551f
c_162 XI5/NET01370 0 0.176433f
c_163 XI5/NET01402 0 0.176433f
c_164 XI5/NET01434 0 0.176433f
c_165 XI5/NET01466 0 0.176433f
c_166 XI5/NET01498 0 0.176433f
c_167 XI5/NET01530 0 0.176433f
c_168 XI5/NET01562 0 0.176433f
c_169 XI5/NET01594 0 0.18066f
c_170 XI5/NET01626 0 0.176433f
c_171 XI5/NET01658 0 0.176433f
c_172 XI5/NET01690 0 0.176433f
c_173 XI5/NET01722 0 0.176433f
c_174 XI5/NET01754 0 0.176433f
c_175 XI5/NET01786 0 0.176433f
c_176 XI5/NET01818 0 0.176433f
c_177 XI5/NET01850 0 0.18066f
c_178 XI5/NET01882 0 0.176433f
c_179 XI5/NET01914 0 0.176433f
c_180 XI5/NET01946 0 0.176433f
c_181 XI5/NET01978 0 0.176433f
c_182 XI5/NET02010 0 0.176433f
c_183 XI5/NET02042 0 0.176433f
c_184 XI5/NET02074 0 0.176433f
c_185 XI5/NET02106 0 0.18066f
c_186 XI5/NET02138 0 0.176433f
c_187 XI5/NET02170 0 0.176433f
c_188 XI5/NET02202 0 0.176433f
c_189 XI5/NET02234 0 0.176433f
c_190 XI5/NET02266 0 0.176433f
c_191 XI5/NET02290 0 0.176433f
c_192 XI5/NET04522 0 0.176433f
c_193 XI5/NET02322 0 0.176433f
c_194 XI5/NET02358 0 0.176433f
c_195 XI5/NET02390 0 0.176433f
c_196 XI5/NET02422 0 0.176433f
c_197 XI5/NET02454 0 0.176433f
c_198 XI5/NET04274 0 0.176433f
c_199 XI5/NET04306 0 0.176433f
c_200 XI5/NET03454 0 0.176433f
c_201 XI5/NET05394 0 0.176433f
c_202 XI5/NET05350 0 0.176433f
c_203 XI5/NET05306 0 0.176433f
c_204 XI5/NET05274 0 0.176433f
c_205 XI5/NET05242 0 0.176433f
c_206 XI5/NET05210 0 0.176433f
c_207 XI5/NET05170 0 0.176433f
c_208 XI5/NET05138 0 0.176433f
c_209 XI5/NET05102 0 0.176433f
c_210 XI5/NET05070 0 0.176433f
c_211 XI5/NET05038 0 0.176433f
c_212 XI5/NET05006 0 0.176433f
c_213 XI5/NET04974 0 0.176433f
c_214 XI5/NET04942 0 0.176433f
c_215 XI5/NET04902 0 0.176433f
c_216 XI5/NET04870 0 0.176433f
c_217 XI5/NET04838 0 0.176433f
c_218 XI5/NET04806 0 0.176433f
c_219 XI5/NET04754 0 0.176433f
c_220 XI5/NET04714 0 0.176433f
c_221 XI5/NET04638 0 0.176433f
c_222 XI5/NET04606 0 0.176433f
c_223 XI5/NET04570 0 0.176433f
c_224 XI5/NET04374 0 0.176433f
c_225 XI5/NET01334 0 0.180551f
c_226 XI5/NET01366 0 0.176433f
c_227 XI5/NET01398 0 0.176433f
c_228 XI5/NET01430 0 0.176433f
c_229 XI5/NET01462 0 0.176433f
c_230 XI5/NET01494 0 0.176433f
c_231 XI5/NET01526 0 0.176433f
c_232 XI5/NET01558 0 0.176433f
c_233 XI5/NET01590 0 0.18066f
c_234 XI5/NET01622 0 0.176433f
c_235 XI5/NET01654 0 0.176433f
c_236 XI5/NET01686 0 0.176433f
c_237 XI5/NET01718 0 0.176433f
c_238 XI5/NET01750 0 0.176433f
c_239 XI5/NET01782 0 0.176433f
c_240 XI5/NET01814 0 0.176433f
c_241 XI5/NET01846 0 0.18066f
c_242 XI5/NET01878 0 0.176433f
c_243 XI5/NET01910 0 0.176433f
c_244 XI5/NET01942 0 0.176433f
c_245 XI5/NET01974 0 0.176433f
c_246 XI5/NET02006 0 0.176433f
c_247 XI5/NET02038 0 0.176433f
c_248 XI5/NET02070 0 0.176433f
c_249 XI5/NET02102 0 0.18066f
c_250 XI5/NET02134 0 0.176433f
c_251 XI5/NET02166 0 0.176433f
c_252 XI5/NET02198 0 0.176433f
c_253 XI5/NET02230 0 0.176433f
c_254 XI5/NET02262 0 0.176433f
c_255 XI5/NET02294 0 0.176433f
c_256 XI5/NET04518 0 0.176433f
c_257 XI5/NET02330 0 0.176433f
c_258 XI5/NET02354 0 0.176433f
c_259 XI5/NET02386 0 0.176433f
c_260 XI5/NET02418 0 0.176433f
c_261 XI5/NET02450 0 0.176433f
c_262 XI5/NET04270 0 0.176433f
c_263 XI5/NET04302 0 0.176433f
c_264 XI5/NET03450 0 0.176433f
c_265 XI5/NET05390 0 0.176433f
c_266 XI5/NET05346 0 0.176433f
c_267 XI5/NET05302 0 0.176433f
c_268 XI5/NET05270 0 0.176433f
c_269 XI5/NET05238 0 0.176433f
c_270 XI5/NET05206 0 0.176433f
c_271 XI5/NET05166 0 0.176433f
c_272 XI5/NET05134 0 0.176433f
c_273 XI5/NET05098 0 0.176433f
c_274 XI5/NET05066 0 0.176433f
c_275 XI5/NET05034 0 0.176433f
c_276 XI5/NET05002 0 0.176433f
c_277 XI5/NET04970 0 0.176433f
c_278 XI5/NET04938 0 0.176433f
c_279 XI5/NET04898 0 0.176433f
c_280 XI5/NET04866 0 0.176433f
c_281 XI5/NET04834 0 0.176433f
c_282 XI5/NET04802 0 0.176433f
c_283 XI5/NET04750 0 0.176433f
c_284 XI5/NET04710 0 0.176433f
c_285 XI5/NET04634 0 0.176433f
c_286 XI5/NET04602 0 0.176433f
c_287 XI5/NET04558 0 0.176433f
c_288 XI5/NET04370 0 0.176433f
c_289 XI5/NET01330 0 0.180551f
c_290 XI5/NET01362 0 0.176433f
c_291 XI5/NET01394 0 0.176433f
c_292 XI5/NET01426 0 0.176433f
c_293 XI5/NET01458 0 0.176433f
c_294 XI5/NET01490 0 0.176433f
c_295 XI5/NET01522 0 0.176433f
c_296 XI5/NET01554 0 0.176433f
c_297 XI5/NET01586 0 0.18066f
c_298 XI5/NET01618 0 0.176433f
c_299 XI5/NET01650 0 0.176433f
c_300 XI5/NET01682 0 0.176433f
c_301 XI5/NET01714 0 0.176433f
c_302 XI5/NET01746 0 0.176433f
c_303 XI5/NET01778 0 0.176433f
c_304 XI5/NET01810 0 0.176433f
c_305 XI5/NET01842 0 0.18066f
c_306 XI5/NET01874 0 0.176433f
c_307 XI5/NET01906 0 0.176433f
c_308 XI5/NET01938 0 0.176433f
c_309 XI5/NET01970 0 0.176433f
c_310 XI5/NET02002 0 0.176433f
c_311 XI5/NET02034 0 0.176433f
c_312 XI5/NET02066 0 0.176433f
c_313 XI5/NET02098 0 0.18066f
c_314 XI5/NET02130 0 0.176433f
c_315 XI5/NET02162 0 0.176433f
c_316 XI5/NET02194 0 0.176433f
c_317 XI5/NET02226 0 0.176433f
c_318 XI5/NET02258 0 0.176433f
c_319 XI5/NET02286 0 0.176433f
c_320 XI5/NET04514 0 0.176433f
c_321 XI5/NET02314 0 0.176433f
c_322 XI5/NET02350 0 0.176433f
c_323 XI5/NET02382 0 0.176433f
c_324 XI5/NET02414 0 0.176433f
c_325 XI5/NET02446 0 0.176433f
c_326 XI5/NET04266 0 0.176433f
c_327 XI5/NET04298 0 0.176433f
c_328 XI5/NET03446 0 0.176433f
c_329 XI5/NET05386 0 0.176433f
c_330 XI5/NET05342 0 0.176433f
c_331 XI5/NET05298 0 0.176433f
c_332 XI5/NET05266 0 0.176433f
c_333 XI5/NET05234 0 0.176433f
c_334 XI5/NET05202 0 0.176433f
c_335 XI5/NET05162 0 0.176433f
c_336 XI5/NET05130 0 0.176433f
c_337 XI5/NET05094 0 0.176433f
c_338 XI5/NET05062 0 0.176433f
c_339 XI5/NET05030 0 0.176433f
c_340 XI5/NET04998 0 0.176433f
c_341 XI5/NET04966 0 0.176433f
c_342 XI5/NET04934 0 0.176433f
c_343 XI5/NET04894 0 0.176433f
c_344 XI5/NET04862 0 0.176433f
c_345 XI5/NET04830 0 0.176433f
c_346 XI5/NET04798 0 0.176433f
c_347 XI5/NET04746 0 0.176433f
c_348 XI5/NET04706 0 0.176433f
c_349 XI5/NET04630 0 0.176433f
c_350 XI5/NET04598 0 0.176433f
c_351 XI5/NET04554 0 0.176433f
c_352 XI5/NET04322 0 0.176433f
c_353 XI5/NET01326 0 0.180551f
c_354 XI5/NET01358 0 0.176433f
c_355 XI5/NET01390 0 0.176433f
c_356 XI5/NET01422 0 0.176433f
c_357 XI5/NET01454 0 0.176433f
c_358 XI5/NET01486 0 0.176433f
c_359 XI5/NET01518 0 0.176433f
c_360 XI5/NET01550 0 0.176433f
c_361 XI5/NET01582 0 0.18066f
c_362 XI5/NET01614 0 0.176433f
c_363 XI5/NET01646 0 0.176433f
c_364 XI5/NET01678 0 0.176433f
c_365 XI5/NET01710 0 0.176433f
c_366 XI5/NET01742 0 0.176433f
c_367 XI5/NET01774 0 0.176433f
c_368 XI5/NET01806 0 0.176433f
c_369 XI5/NET01838 0 0.18066f
c_370 XI5/NET01870 0 0.176433f
c_371 XI5/NET01902 0 0.176433f
c_372 XI5/NET01934 0 0.176433f
c_373 XI5/NET01966 0 0.176433f
c_374 XI5/NET01998 0 0.176433f
c_375 XI5/NET02030 0 0.176433f
c_376 XI5/NET02062 0 0.176433f
c_377 XI5/NET02094 0 0.18066f
c_378 XI5/NET02126 0 0.176433f
c_379 XI5/NET02158 0 0.176433f
c_380 XI5/NET02190 0 0.176433f
c_381 XI5/NET02222 0 0.176433f
c_382 XI5/NET02254 0 0.176433f
c_383 XI5/NET02306 0 0.176433f
c_384 XI5/NET04510 0 0.176433f
c_385 XI5/NET02318 0 0.176433f
c_386 XI5/NET02346 0 0.176433f
c_387 XI5/NET02378 0 0.176433f
c_388 XI5/NET02410 0 0.176433f
c_389 XI5/NET02442 0 0.176433f
c_390 XI5/NET04262 0 0.176433f
c_391 XI5/NET04294 0 0.176433f
c_392 XI5/NET03442 0 0.176433f
c_393 XI5/NET05382 0 0.176433f
c_394 XI5/NET05338 0 0.176433f
c_395 XI5/NET05294 0 0.176433f
c_396 XI5/NET05262 0 0.176433f
c_397 XI5/NET05230 0 0.176433f
c_398 XI5/NET05198 0 0.176433f
c_399 XI5/NET05158 0 0.176433f
c_400 XI5/NET05126 0 0.176433f
c_401 XI5/NET05090 0 0.176433f
c_402 XI5/NET05058 0 0.176433f
c_403 XI5/NET05026 0 0.176433f
c_404 XI5/NET04994 0 0.176433f
c_405 XI5/NET04962 0 0.176433f
c_406 XI5/NET04930 0 0.176433f
c_407 XI5/NET04890 0 0.176433f
c_408 XI5/NET04858 0 0.176433f
c_409 XI5/NET04826 0 0.176433f
c_410 XI5/NET04794 0 0.176433f
c_411 XI5/NET04742 0 0.176433f
c_412 XI5/NET04694 0 0.176433f
c_413 XI5/NET04626 0 0.176433f
c_414 XI5/NET04594 0 0.176433f
c_415 XI5/NET04550 0 0.176433f
c_416 XI5/NET03002 0 0.176433f
c_417 XI5/NET01322 0 0.180551f
c_418 XI5/NET01354 0 0.176433f
c_419 XI5/NET01386 0 0.176433f
c_420 XI5/NET01418 0 0.176433f
c_421 XI5/NET01450 0 0.176433f
c_422 XI5/NET01482 0 0.176433f
c_423 XI5/NET01514 0 0.176433f
c_424 XI5/NET01546 0 0.176433f
c_425 XI5/NET01578 0 0.18066f
c_426 XI5/NET01610 0 0.176433f
c_427 XI5/NET01642 0 0.176433f
c_428 XI5/NET01674 0 0.176433f
c_429 XI5/NET01706 0 0.176433f
c_430 XI5/NET01738 0 0.176433f
c_431 XI5/NET01770 0 0.176433f
c_432 XI5/NET01802 0 0.176433f
c_433 XI5/NET01834 0 0.18066f
c_434 XI5/NET01866 0 0.176433f
c_435 XI5/NET01898 0 0.176433f
c_436 XI5/NET01930 0 0.176433f
c_437 XI5/NET01962 0 0.176433f
c_438 XI5/NET01994 0 0.176433f
c_439 XI5/NET02026 0 0.176433f
c_440 XI5/NET02058 0 0.176433f
c_441 XI5/NET02090 0 0.18066f
c_442 XI5/NET02122 0 0.176433f
c_443 XI5/NET02154 0 0.176433f
c_444 XI5/NET02186 0 0.176433f
c_445 XI5/NET02218 0 0.176433f
c_446 XI5/NET02250 0 0.176433f
c_447 XI5/NET02298 0 0.176433f
c_448 XI5/NET04434 0 0.176433f
c_449 XI5/NET02334 0 0.176433f
c_450 XI5/NET02342 0 0.176433f
c_451 XI5/NET02374 0 0.176433f
c_452 XI5/NET02406 0 0.176433f
c_453 XI5/NET02438 0 0.176433f
c_454 XI5/NET04258 0 0.176433f
c_455 XI5/NET04290 0 0.176433f
c_456 XI5/NET03438 0 0.176433f
c_457 XI5/NET05378 0 0.176433f
c_458 XI5/NET05334 0 0.176433f
c_459 XI5/NET05290 0 0.176433f
c_460 XI5/NET05258 0 0.176433f
c_461 XI5/NET05226 0 0.176433f
c_462 XI5/NET05194 0 0.176433f
c_463 XI5/NET05154 0 0.176433f
c_464 XI5/NET05122 0 0.176433f
c_465 XI5/NET05086 0 0.176433f
c_466 XI5/NET05054 0 0.176433f
c_467 XI5/NET05022 0 0.176433f
c_468 XI5/NET04990 0 0.176433f
c_469 XI5/NET04958 0 0.176433f
c_470 XI5/NET04926 0 0.176433f
c_471 XI5/NET04886 0 0.176433f
c_472 XI5/NET04854 0 0.176433f
c_473 XI5/NET04822 0 0.176433f
c_474 XI5/NET04790 0 0.176433f
c_475 XI5/NET04738 0 0.176433f
c_476 XI5/NET04666 0 0.176433f
c_477 XI5/NET04622 0 0.176433f
c_478 XI5/NET04590 0 0.176433f
c_479 XI5/NET04546 0 0.176433f
c_480 XI5/NET02746 0 0.176433f
c_481 XI5/NET01318 0 0.138298f
c_482 XI5/NET01350 0 0.136314f
c_483 XI5/NET01382 0 0.136314f
c_484 XI5/NET01414 0 0.136314f
c_485 XI5/NET01446 0 0.136314f
c_486 XI5/NET01478 0 0.136314f
c_487 XI5/NET01510 0 0.136314f
c_488 XI5/NET01542 0 0.136314f
c_489 XI5/NET01574 0 0.138908f
c_490 XI5/NET01606 0 0.136314f
c_491 XI5/NET01638 0 0.136314f
c_492 XI5/NET01670 0 0.136314f
c_493 XI5/NET01702 0 0.136314f
c_494 XI5/NET01734 0 0.136314f
c_495 XI5/NET01766 0 0.136314f
c_496 XI5/NET01798 0 0.136314f
c_497 XI5/NET01830 0 0.138908f
c_498 XI5/NET01862 0 0.136314f
c_499 XI5/NET01894 0 0.136314f
c_500 XI5/NET01926 0 0.136314f
c_501 XI5/NET01958 0 0.136314f
c_502 XI5/NET01990 0 0.136314f
c_503 XI5/NET02022 0 0.136314f
c_504 XI5/NET02054 0 0.136314f
c_505 XI5/NET02086 0 0.138908f
c_506 XI5/NET02118 0 0.136314f
c_507 XI5/NET02150 0 0.136314f
c_508 XI5/NET02182 0 0.136314f
c_509 XI5/NET02214 0 0.136314f
c_510 XI5/NET02246 0 0.136314f
c_511 XI5/NET02302 0 0.136314f
c_512 XI5/NET04394 0 0.136314f
*
.include "ROM_MACRO.pex.spi.ROM_MACRO.pxi"
*
.ends
*
*
